
module fpu_DW01_inc_0 ( A, SUM );
  input [21:0] A;
  output [21:0] SUM;

  wire   [21:2] carry;

  HADDX1_RVT U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1_RVT U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1_RVT U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1_RVT U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1_RVT U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1_RVT U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1_RVT U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1_RVT U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1_RVT U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1_RVT U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1_RVT U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1_RVT U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1_RVT U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[21]), .A2(A[21]), .Y(SUM[21]) );
endmodule


module fpu_DW01_inc_1 ( A, SUM );
  input [21:0] A;
  output [21:0] SUM;

  wire   [21:2] carry;

  HADDX1_RVT U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1_RVT U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1_RVT U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1_RVT U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1_RVT U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1_RVT U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1_RVT U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1_RVT U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1_RVT U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1_RVT U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1_RVT U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1_RVT U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1_RVT U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[21]), .A2(A[21]), .Y(SUM[21]) );
endmodule


module fpu_DW01_inc_2 ( A, SUM );
  input [9:0] A;
  output [9:0] SUM;
  wire   n1;
  wire   [9:2] carry;

  HADDX1_RVT U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(n1), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  INVX1_RVT U2 ( .A(SUM[0]), .Y(n1) );
  XOR2X1_RVT U3 ( .A1(carry[9]), .A2(A[9]), .Y(SUM[9]) );
endmodule


module fpu_DW01_add_2 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;

  wire   [8:1] carry;

  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(SUM[8]), .S(SUM[7])
         );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module fpu_DW01_inc_3 ( A, SUM );
  input [21:0] A;
  output [21:0] SUM;

  wire   [21:2] carry;

  HADDX1_RVT U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1_RVT U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1_RVT U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1_RVT U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1_RVT U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1_RVT U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1_RVT U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1_RVT U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1_RVT U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1_RVT U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1_RVT U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1_RVT U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1_RVT U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[21]), .A2(A[21]), .Y(SUM[21]) );
endmodule


module fpu_DW01_inc_4 ( A, SUM );
  input [21:0] A;
  output [21:0] SUM;

  wire   [21:2] carry;

  HADDX1_RVT U1_1_20 ( .A0(A[20]), .B0(carry[20]), .C1(carry[21]), .SO(SUM[20]) );
  HADDX1_RVT U1_1_19 ( .A0(A[19]), .B0(carry[19]), .C1(carry[20]), .SO(SUM[19]) );
  HADDX1_RVT U1_1_18 ( .A0(A[18]), .B0(carry[18]), .C1(carry[19]), .SO(SUM[18]) );
  HADDX1_RVT U1_1_17 ( .A0(A[17]), .B0(carry[17]), .C1(carry[18]), .SO(SUM[17]) );
  HADDX1_RVT U1_1_16 ( .A0(A[16]), .B0(carry[16]), .C1(carry[17]), .SO(SUM[16]) );
  HADDX1_RVT U1_1_15 ( .A0(A[15]), .B0(carry[15]), .C1(carry[16]), .SO(SUM[15]) );
  HADDX1_RVT U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1_RVT U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1_RVT U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1_RVT U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1_RVT U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1_RVT U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1_RVT U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1_RVT U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[21]), .A2(A[21]), .Y(SUM[21]) );
endmodule


module fpu_DW01_inc_5 ( A, SUM );
  input [7:0] A;
  output [7:0] SUM;

  wire   [7:2] carry;

  HADDX1_RVT U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1_RVT U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1_RVT U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1_RVT U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1_RVT U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1_RVT U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX1_RVT U1 ( .A(A[0]), .Y(SUM[0]) );
  XOR2X1_RVT U2 ( .A1(carry[7]), .A2(A[7]), .Y(SUM[7]) );
endmodule


module fpu_DW01_inc_6 ( A, SUM );
  input [47:0] A;
  output [47:0] SUM;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [47:2] carry;

  HADDX1_RVT U1_1_46 ( .A0(A[46]), .B0(carry[46]), .C1(carry[47]), .SO(SUM[46]) );
  HADDX1_RVT U1_1_45 ( .A0(A[45]), .B0(carry[45]), .C1(carry[46]), .SO(SUM[45]) );
  HADDX1_RVT U1_1_44 ( .A0(A[44]), .B0(carry[44]), .C1(carry[45]), .SO(SUM[44]) );
  HADDX1_RVT U1_1_43 ( .A0(A[43]), .B0(carry[43]), .C1(carry[44]), .SO(SUM[43]) );
  HADDX1_RVT U1_1_42 ( .A0(A[42]), .B0(carry[42]), .C1(carry[43]), .SO(SUM[42]) );
  HADDX1_RVT U1_1_41 ( .A0(A[41]), .B0(carry[41]), .C1(carry[42]), .SO(SUM[41]) );
  HADDX1_RVT U1_1_40 ( .A0(A[40]), .B0(carry[40]), .C1(carry[41]), .SO(SUM[40]) );
  HADDX1_RVT U1_1_39 ( .A0(A[39]), .B0(carry[39]), .C1(carry[40]), .SO(SUM[39]) );
  HADDX1_RVT U1_1_38 ( .A0(A[38]), .B0(carry[38]), .C1(carry[39]), .SO(SUM[38]) );
  HADDX1_RVT U1_1_37 ( .A0(A[37]), .B0(carry[37]), .C1(carry[38]), .SO(SUM[37]) );
  HADDX1_RVT U1_1_36 ( .A0(A[36]), .B0(carry[36]), .C1(carry[37]), .SO(SUM[36]) );
  HADDX1_RVT U1_1_35 ( .A0(A[35]), .B0(carry[35]), .C1(carry[36]), .SO(SUM[35]) );
  HADDX1_RVT U1_1_34 ( .A0(A[34]), .B0(carry[34]), .C1(carry[35]), .SO(SUM[34]) );
  HADDX1_RVT U1_1_33 ( .A0(A[33]), .B0(carry[33]), .C1(carry[34]), .SO(SUM[33]) );
  HADDX1_RVT U1_1_32 ( .A0(A[32]), .B0(carry[32]), .C1(carry[33]), .SO(SUM[32]) );
  HADDX1_RVT U1_1_31 ( .A0(A[31]), .B0(carry[31]), .C1(carry[32]), .SO(SUM[31]) );
  HADDX1_RVT U1_1_30 ( .A0(A[30]), .B0(carry[30]), .C1(carry[31]), .SO(SUM[30]) );
  HADDX1_RVT U1_1_29 ( .A0(A[29]), .B0(carry[29]), .C1(carry[30]), .SO(SUM[29]) );
  HADDX1_RVT U1_1_28 ( .A0(A[28]), .B0(carry[28]), .C1(carry[29]), .SO(SUM[28]) );
  HADDX1_RVT U1_1_27 ( .A0(A[27]), .B0(carry[27]), .C1(carry[28]), .SO(SUM[27]) );
  HADDX1_RVT U1_1_26 ( .A0(A[26]), .B0(carry[26]), .C1(carry[27]), .SO(SUM[26]) );
  HADDX1_RVT U1_1_25 ( .A0(A[25]), .B0(carry[25]), .C1(carry[26]), .SO(SUM[25]) );
  HADDX1_RVT U1_1_24 ( .A0(A[24]), .B0(carry[24]), .C1(carry[25]), .SO(SUM[24]) );
  NOR4X0_RVT U1 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .Y(carry[24]) );
  NAND4X0_RVT U2 ( .A1(A[8]), .A2(A[7]), .A3(A[9]), .A4(n5), .Y(n4) );
  AND3X1_RVT U3 ( .A1(A[5]), .A2(A[4]), .A3(A[6]), .Y(n5) );
  NAND4X0_RVT U4 ( .A1(A[2]), .A2(A[23]), .A3(A[3]), .A4(n6), .Y(n3) );
  AND3X1_RVT U5 ( .A1(A[21]), .A2(A[20]), .A3(A[22]), .Y(n6) );
  NAND4X0_RVT U6 ( .A1(A[19]), .A2(A[18]), .A3(A[1]), .A4(n7), .Y(n2) );
  AND3X1_RVT U7 ( .A1(A[16]), .A2(A[15]), .A3(A[17]), .Y(n7) );
  NAND4X0_RVT U8 ( .A1(A[13]), .A2(A[12]), .A3(A[14]), .A4(n8), .Y(n1) );
  AND3X1_RVT U9 ( .A1(A[10]), .A2(A[0]), .A3(A[11]), .Y(n8) );
  XOR2X1_RVT U10 ( .A1(carry[47]), .A2(A[47]), .Y(SUM[47]) );
endmodule


module fpu_DW01_sub_24 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [25:0] carry;

  FADDX1_RVT U2_22 ( .A(A[22]), .B(n23), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1_RVT U2_21 ( .A(A[21]), .B(n22), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1_RVT U2_20 ( .A(A[20]), .B(n21), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1_RVT U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1_RVT U2_12 ( .A(A[12]), .B(n13), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1_RVT U2_10 ( .A(A[10]), .B(n11), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1_RVT U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n4), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_13 ( .A(A[13]), .B(n14), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1_RVT U2_11 ( .A(A[11]), .B(n12), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1_RVT U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1_RVT U2_15 ( .A(A[15]), .B(n16), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n6), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1_RVT U2_9 ( .A(A[9]), .B(n10), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n2), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FADDX1_RVT U2_18 ( .A(A[18]), .B(n19), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1_RVT U2_19 ( .A(A[19]), .B(n20), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1_RVT U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1_RVT U2_17 ( .A(A[17]), .B(n18), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1_RVT U2_7 ( .A(A[7]), .B(n8), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1_RVT U2_23 ( .A(A[23]), .B(n24), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n3), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INVX0_RVT U1 ( .A(B[2]), .Y(n3) );
  INVX0_RVT U2 ( .A(B[23]), .Y(n24) );
  INVX0_RVT U3 ( .A(B[21]), .Y(n22) );
  INVX0_RVT U4 ( .A(B[22]), .Y(n23) );
  INVX0_RVT U5 ( .A(B[20]), .Y(n21) );
  INVX0_RVT U6 ( .A(B[1]), .Y(n2) );
  XNOR2X1_RVT U7 ( .A1(A[0]), .A2(n1), .Y(DIFF[0]) );
  INVX1_RVT U8 ( .A(carry[24]), .Y(DIFF[24]) );
  INVX1_RVT U9 ( .A(B[7]), .Y(n8) );
  INVX1_RVT U10 ( .A(B[17]), .Y(n18) );
  INVX1_RVT U11 ( .A(B[8]), .Y(n9) );
  INVX1_RVT U12 ( .A(B[19]), .Y(n20) );
  INVX1_RVT U13 ( .A(B[18]), .Y(n19) );
  INVX1_RVT U14 ( .A(B[0]), .Y(n1) );
  OR2X1_RVT U15 ( .A1(n1), .A2(A[0]), .Y(carry[1]) );
  INVX1_RVT U16 ( .A(B[9]), .Y(n10) );
  INVX1_RVT U17 ( .A(B[5]), .Y(n6) );
  INVX1_RVT U18 ( .A(B[15]), .Y(n16) );
  INVX1_RVT U19 ( .A(B[4]), .Y(n5) );
  INVX1_RVT U20 ( .A(B[6]), .Y(n7) );
  INVX1_RVT U21 ( .A(B[11]), .Y(n12) );
  INVX1_RVT U22 ( .A(B[13]), .Y(n14) );
  INVX1_RVT U23 ( .A(B[3]), .Y(n4) );
  INVX1_RVT U24 ( .A(B[16]), .Y(n17) );
  INVX1_RVT U25 ( .A(B[10]), .Y(n11) );
  INVX1_RVT U26 ( .A(B[12]), .Y(n13) );
  INVX1_RVT U27 ( .A(B[14]), .Y(n15) );
endmodule


module fpu_DW01_sub_25 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24;
  wire   [25:0] carry;

  FADDX1_RVT U2_22 ( .A(A[22]), .B(n23), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1_RVT U2_21 ( .A(A[21]), .B(n22), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1_RVT U2_20 ( .A(A[20]), .B(n21), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1_RVT U2_18 ( .A(A[18]), .B(n19), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1_RVT U2_19 ( .A(A[19]), .B(n20), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1_RVT U2_17 ( .A(A[17]), .B(n18), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1_RVT U2_15 ( .A(A[15]), .B(n16), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1_RVT U2_16 ( .A(A[16]), .B(n17), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1_RVT U2_14 ( .A(A[14]), .B(n15), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1_RVT U2_13 ( .A(A[13]), .B(n14), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1_RVT U2_12 ( .A(A[12]), .B(n13), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1_RVT U2_11 ( .A(A[11]), .B(n12), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1_RVT U2_10 ( .A(A[10]), .B(n11), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1_RVT U2_9 ( .A(A[9]), .B(n10), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  FADDX1_RVT U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1_RVT U2_7 ( .A(A[7]), .B(n8), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n2), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FADDX1_RVT U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n4), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n6), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n7), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1_RVT U2_23 ( .A(A[23]), .B(n24), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n3), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  INVX0_RVT U1 ( .A(B[2]), .Y(n3) );
  INVX0_RVT U2 ( .A(B[5]), .Y(n6) );
  INVX0_RVT U3 ( .A(B[6]), .Y(n7) );
  INVX0_RVT U4 ( .A(B[3]), .Y(n4) );
  INVX0_RVT U5 ( .A(B[12]), .Y(n13) );
  INVX0_RVT U6 ( .A(B[13]), .Y(n14) );
  INVX0_RVT U7 ( .A(B[11]), .Y(n12) );
  INVX0_RVT U8 ( .A(B[23]), .Y(n24) );
  INVX0_RVT U9 ( .A(B[14]), .Y(n15) );
  INVX1_RVT U10 ( .A(carry[24]), .Y(DIFF[24]) );
  INVX1_RVT U11 ( .A(B[0]), .Y(n1) );
  XNOR2X1_RVT U12 ( .A1(A[0]), .A2(n1), .Y(DIFF[0]) );
  INVX1_RVT U13 ( .A(B[4]), .Y(n5) );
  INVX1_RVT U14 ( .A(B[1]), .Y(n2) );
  OR2X1_RVT U15 ( .A1(n1), .A2(A[0]), .Y(carry[1]) );
  INVX1_RVT U16 ( .A(B[7]), .Y(n8) );
  INVX1_RVT U17 ( .A(B[8]), .Y(n9) );
  INVX1_RVT U18 ( .A(B[9]), .Y(n10) );
  INVX1_RVT U19 ( .A(B[10]), .Y(n11) );
  INVX1_RVT U20 ( .A(B[16]), .Y(n17) );
  INVX1_RVT U21 ( .A(B[15]), .Y(n16) );
  INVX1_RVT U22 ( .A(B[17]), .Y(n18) );
  INVX1_RVT U23 ( .A(B[19]), .Y(n20) );
  INVX1_RVT U24 ( .A(B[18]), .Y(n19) );
  INVX1_RVT U25 ( .A(B[20]), .Y(n21) );
  INVX1_RVT U26 ( .A(B[21]), .Y(n22) );
  INVX1_RVT U27 ( .A(B[22]), .Y(n23) );
endmodule


module fpu_DW01_sub_26 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [25:0] carry;

  FADDX1_RVT U2_4 ( .A(A[4]), .B(n14), .CI(carry[4]), .CO(carry[5]), .S(
        DIFF[4]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n16), .CI(carry[6]), .CO(carry[7]), .S(
        DIFF[6]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n15), .CI(carry[5]), .CO(carry[6]), .S(
        DIFF[5]) );
  FADDX1_RVT U2_9 ( .A(A[9]), .B(n19), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  FADDX1_RVT U2_16 ( .A(A[16]), .B(n20), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1_RVT U2_18 ( .A(A[18]), .B(n22), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1_RVT U2_17 ( .A(A[17]), .B(n21), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1_RVT U2_19 ( .A(A[19]), .B(n23), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1_RVT U2_20 ( .A(A[20]), .B(n10), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1_RVT U2_23 ( .A(A[23]), .B(n13), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1_RVT U2_21 ( .A(A[21]), .B(n11), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1_RVT U2_22 ( .A(A[22]), .B(n12), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1_RVT U2_15 ( .A(A[15]), .B(n9), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1_RVT U2_14 ( .A(A[14]), .B(n8), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1_RVT U2_7 ( .A(A[7]), .B(n17), .CI(carry[7]), .CO(carry[8]), .S(
        DIFF[7]) );
  FADDX1_RVT U2_10 ( .A(A[10]), .B(n4), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1_RVT U2_12 ( .A(A[12]), .B(n6), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1_RVT U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1_RVT U2_13 ( .A(A[13]), .B(n7), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n25), .CI(carry[2]), .CO(carry[3]), .S(
        DIFF[2]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n2), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_8 ( .A(A[8]), .B(n18), .CI(carry[8]), .CO(carry[9]), .S(
        DIFF[8]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n24), .CI(carry[1]), .CO(carry[2]), .S(
        DIFF[1]) );
  INVX1_RVT U1 ( .A(B[6]), .Y(n16) );
  OR2X1_RVT U2 ( .A1(n3), .A2(A[0]), .Y(carry[1]) );
  INVX1_RVT U3 ( .A(B[8]), .Y(n18) );
  INVX1_RVT U4 ( .A(B[5]), .Y(n15) );
  INVX1_RVT U5 ( .A(B[2]), .Y(n25) );
  INVX1_RVT U6 ( .A(B[12]), .Y(n6) );
  INVX1_RVT U7 ( .A(B[7]), .Y(n17) );
  INVX1_RVT U8 ( .A(B[20]), .Y(n10) );
  INVX1_RVT U9 ( .A(B[11]), .Y(n5) );
  INVX1_RVT U10 ( .A(B[10]), .Y(n4) );
  INVX1_RVT U11 ( .A(B[9]), .Y(n19) );
  INVX1_RVT U12 ( .A(B[13]), .Y(n7) );
  INVX1_RVT U13 ( .A(B[14]), .Y(n8) );
  INVX1_RVT U14 ( .A(B[15]), .Y(n9) );
  INVX1_RVT U15 ( .A(B[0]), .Y(n3) );
  INVX1_RVT U16 ( .A(B[21]), .Y(n11) );
  INVX1_RVT U17 ( .A(B[3]), .Y(n2) );
  INVX1_RVT U18 ( .A(B[1]), .Y(n24) );
  XNOR2X1_RVT U19 ( .A1(A[0]), .A2(n3), .Y(DIFF[0]) );
  INVX1_RVT U20 ( .A(B[4]), .Y(n14) );
  INVX0_RVT U21 ( .A(B[22]), .Y(n12) );
  INVX1_RVT U22 ( .A(B[23]), .Y(n13) );
  INVX0_RVT U23 ( .A(B[19]), .Y(n23) );
  INVX0_RVT U24 ( .A(B[17]), .Y(n21) );
  INVX1_RVT U25 ( .A(B[18]), .Y(n22) );
  INVX0_RVT U26 ( .A(B[16]), .Y(n20) );
  INVX1_RVT U27 ( .A(carry[24]), .Y(DIFF[24]) );
endmodule


module fpu_DW01_sub_27 ( A, B, CI, DIFF, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [25:0] carry;

  FADDX1_RVT U2_4 ( .A(A[4]), .B(n14), .CI(carry[4]), .CO(carry[5]), .S(
        DIFF[4]) );
  FADDX1_RVT U2_8 ( .A(A[8]), .B(n18), .CI(carry[8]), .CO(carry[9]), .S(
        DIFF[8]) );
  FADDX1_RVT U2_9 ( .A(A[9]), .B(n19), .CI(carry[9]), .CO(carry[10]), .S(
        DIFF[9]) );
  FADDX1_RVT U2_7 ( .A(A[7]), .B(n17), .CI(carry[7]), .CO(carry[8]), .S(
        DIFF[7]) );
  FADDX1_RVT U2_20 ( .A(A[20]), .B(n10), .CI(carry[20]), .CO(carry[21]), .S(
        DIFF[20]) );
  FADDX1_RVT U2_18 ( .A(A[18]), .B(n22), .CI(carry[18]), .CO(carry[19]), .S(
        DIFF[18]) );
  FADDX1_RVT U2_19 ( .A(A[19]), .B(n23), .CI(carry[19]), .CO(carry[20]), .S(
        DIFF[19]) );
  FADDX1_RVT U2_22 ( .A(A[22]), .B(n12), .CI(carry[22]), .CO(carry[23]), .S(
        DIFF[22]) );
  FADDX1_RVT U2_21 ( .A(A[21]), .B(n11), .CI(carry[21]), .CO(carry[22]), .S(
        DIFF[21]) );
  FADDX1_RVT U2_17 ( .A(A[17]), .B(n21), .CI(carry[17]), .CO(carry[18]), .S(
        DIFF[17]) );
  FADDX1_RVT U2_16 ( .A(A[16]), .B(n20), .CI(carry[16]), .CO(carry[17]), .S(
        DIFF[16]) );
  FADDX1_RVT U2_15 ( .A(A[15]), .B(n9), .CI(carry[15]), .CO(carry[16]), .S(
        DIFF[15]) );
  FADDX1_RVT U2_14 ( .A(A[14]), .B(n8), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1_RVT U2_10 ( .A(A[10]), .B(n4), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1_RVT U2_12 ( .A(A[12]), .B(n6), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1_RVT U2_11 ( .A(A[11]), .B(n5), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1_RVT U2_13 ( .A(A[13]), .B(n7), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n2), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n16), .CI(carry[6]), .CO(carry[7]), .S(
        DIFF[6]) );
  FADDX1_RVT U2_23 ( .A(A[23]), .B(n13), .CI(carry[23]), .CO(carry[24]), .S(
        DIFF[23]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n25), .CI(carry[2]), .CO(carry[3]), .S(
        DIFF[2]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n15), .CI(carry[5]), .CO(carry[6]), .S(
        DIFF[5]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n24), .CI(carry[1]), .CO(carry[2]), .S(
        DIFF[1]) );
  INVX1_RVT U1 ( .A(B[6]), .Y(n16) );
  INVX1_RVT U2 ( .A(B[8]), .Y(n18) );
  INVX1_RVT U3 ( .A(B[5]), .Y(n15) );
  INVX1_RVT U4 ( .A(B[2]), .Y(n25) );
  INVX1_RVT U5 ( .A(B[7]), .Y(n17) );
  INVX1_RVT U6 ( .A(B[10]), .Y(n4) );
  INVX1_RVT U7 ( .A(B[4]), .Y(n14) );
  INVX1_RVT U8 ( .A(B[9]), .Y(n19) );
  INVX1_RVT U9 ( .A(B[13]), .Y(n7) );
  OR2X2_RVT U10 ( .A1(n3), .A2(A[0]), .Y(carry[1]) );
  INVX1_RVT U11 ( .A(B[0]), .Y(n3) );
  INVX1_RVT U12 ( .A(B[1]), .Y(n24) );
  INVX1_RVT U13 ( .A(B[11]), .Y(n5) );
  INVX1_RVT U14 ( .A(B[3]), .Y(n2) );
  INVX1_RVT U15 ( .A(B[14]), .Y(n8) );
  XNOR2X1_RVT U16 ( .A1(A[0]), .A2(n3), .Y(DIFF[0]) );
  INVX1_RVT U17 ( .A(carry[24]), .Y(DIFF[24]) );
  INVX1_RVT U18 ( .A(B[23]), .Y(n13) );
  INVX0_RVT U19 ( .A(B[12]), .Y(n6) );
  INVX1_RVT U20 ( .A(B[15]), .Y(n9) );
  INVX0_RVT U21 ( .A(B[16]), .Y(n20) );
  INVX1_RVT U22 ( .A(B[17]), .Y(n21) );
  INVX1_RVT U23 ( .A(B[21]), .Y(n11) );
  INVX1_RVT U24 ( .A(B[22]), .Y(n12) );
  INVX1_RVT U25 ( .A(B[19]), .Y(n23) );
  INVX0_RVT U26 ( .A(B[18]), .Y(n22) );
  INVX1_RVT U27 ( .A(B[20]), .Y(n10) );
endmodule


module fpu_DW01_add_3 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;

  wire   [24:1] carry;

  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  XOR2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
  AND2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
endmodule


module fpu_DW01_add_4 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;

  wire   [24:1] carry;

  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  AND2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
  XOR2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
endmodule


module fpu_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101;

  AND2X1_RVT U3 ( .A1(n54), .A2(n14), .Y(n20) );
  AOI21X1_RVT U4 ( .A1(n52), .A2(n53), .A3(SH[7]), .Y(B[3]) );
  MUX21X1_RVT U5 ( .A1(n57), .A2(n58), .S0(n15), .Y(n52) );
  INVX0_RVT U6 ( .A(n6), .Y(n11) );
  INVX0_RVT U7 ( .A(n4), .Y(n10) );
  AND2X1_RVT U8 ( .A1(SH[0]), .A2(n18), .Y(n7) );
  AND2X1_RVT U9 ( .A1(n59), .A2(n79), .Y(n1) );
  INVX1_RVT U10 ( .A(n51), .Y(n15) );
  INVX1_RVT U11 ( .A(n89), .Y(n16) );
  AND2X1_RVT U12 ( .A1(n19), .A2(SH[1]), .Y(n2) );
  INVX1_RVT U13 ( .A(n3), .Y(n13) );
  INVX1_RVT U14 ( .A(n3), .Y(n12) );
  NAND2X0_RVT U15 ( .A1(n19), .A2(n18), .Y(n3) );
  INVX1_RVT U16 ( .A(n5), .Y(n8) );
  AO221X1_RVT U17 ( .A1(n20), .A2(n47), .A3(n1), .A4(n25), .A5(n48), .Y(B[4])
         );
  INVX1_RVT U18 ( .A(n4), .Y(n9) );
  NAND2X0_RVT U19 ( .A1(SH[0]), .A2(SH[1]), .Y(n4) );
  INVX1_RVT U20 ( .A(SH[0]), .Y(n19) );
  INVX1_RVT U21 ( .A(SH[1]), .Y(n18) );
  INVX1_RVT U22 ( .A(SH[2]), .Y(n17) );
  NAND2X0_RVT U23 ( .A1(SH[0]), .A2(n18), .Y(n5) );
  INVX1_RVT U24 ( .A(SH[7]), .Y(n14) );
  NAND2X0_RVT U25 ( .A1(n19), .A2(SH[1]), .Y(n6) );
  AO222X1_RVT U26 ( .A1(n20), .A2(n21), .A3(n22), .A4(n23), .A5(n1), .A6(n24), 
        .Y(B[9]) );
  AO222X1_RVT U27 ( .A1(n20), .A2(n25), .A3(n22), .A4(n26), .A5(n1), .A6(n27), 
        .Y(B[8]) );
  AO221X1_RVT U28 ( .A1(n20), .A2(n28), .A3(n1), .A4(n29), .A5(n30), .Y(B[7])
         );
  AO222X1_RVT U29 ( .A1(n31), .A2(n32), .A3(n33), .A4(n34), .A5(n35), .A6(n36), 
        .Y(n30) );
  AO221X1_RVT U30 ( .A1(n20), .A2(n37), .A3(n1), .A4(n38), .A5(n39), .Y(B[6])
         );
  AO222X1_RVT U31 ( .A1(n35), .A2(n40), .A3(n33), .A4(n41), .A5(n31), .A6(n42), 
        .Y(n39) );
  AO221X1_RVT U32 ( .A1(n20), .A2(n43), .A3(n1), .A4(n21), .A5(n44), .Y(B[5])
         );
  AO222X1_RVT U33 ( .A1(n35), .A2(n24), .A3(n33), .A4(n45), .A5(n31), .A6(n46), 
        .Y(n44) );
  AO222X1_RVT U34 ( .A1(n35), .A2(n27), .A3(n33), .A4(n49), .A5(n31), .A6(n50), 
        .Y(n48) );
  AND4X1_RVT U35 ( .A1(n16), .A2(n17), .A3(n51), .A4(n14), .Y(n31) );
  AND2X1_RVT U36 ( .A1(n22), .A2(SH[2]), .Y(n33) );
  NAND2X0_RVT U37 ( .A1(n54), .A2(n55), .Y(n53) );
  AO221X1_RVT U38 ( .A1(A[4]), .A2(n7), .A3(A[3]), .A4(n12), .A5(n56), .Y(n55)
         );
  AO22X1_RVT U39 ( .A1(A[5]), .A2(n2), .A3(A[6]), .A4(n9), .Y(n56) );
  AOI222X1_RVT U40 ( .A1(n28), .A2(n59), .A3(n29), .A4(n60), .A5(n36), .A6(n61), .Y(n58) );
  AO221X1_RVT U41 ( .A1(A[8]), .A2(n7), .A3(A[7]), .A4(n13), .A5(n62), .Y(n28)
         );
  AO22X1_RVT U42 ( .A1(A[9]), .A2(n11), .A3(A[10]), .A4(n10), .Y(n62) );
  NAND2X0_RVT U43 ( .A1(n16), .A2(n63), .Y(n57) );
  OA21X1_RVT U44 ( .A1(n64), .A2(n65), .A3(n14), .Y(B[2]) );
  MUX21X1_RVT U45 ( .A1(n66), .A2(n67), .S0(n15), .Y(n65) );
  AO222X1_RVT U46 ( .A1(n61), .A2(n40), .A3(n60), .A4(n38), .A5(n59), .A6(n37), 
        .Y(n67) );
  AO221X1_RVT U47 ( .A1(A[7]), .A2(n7), .A3(A[6]), .A4(n13), .A5(n68), .Y(n37)
         );
  AO22X1_RVT U48 ( .A1(A[8]), .A2(n2), .A3(A[9]), .A4(n9), .Y(n68) );
  OA21X1_RVT U49 ( .A1(n69), .A2(n70), .A3(n54), .Y(n64) );
  AO22X1_RVT U50 ( .A1(A[2]), .A2(n13), .A3(A[3]), .A4(n7), .Y(n70) );
  AO22X1_RVT U51 ( .A1(A[4]), .A2(n2), .A3(A[5]), .A4(n9), .Y(n69) );
  AND2X1_RVT U52 ( .A1(n32), .A2(n20), .Y(B[23]) );
  AND2X1_RVT U53 ( .A1(n20), .A2(n42), .Y(B[22]) );
  AND2X1_RVT U54 ( .A1(n20), .A2(n46), .Y(B[21]) );
  AND2X1_RVT U55 ( .A1(n20), .A2(n50), .Y(B[20]) );
  OA21X1_RVT U56 ( .A1(n71), .A2(n72), .A3(n14), .Y(B[1]) );
  MUX21X1_RVT U57 ( .A1(n73), .A2(n74), .S0(n15), .Y(n72) );
  AO222X1_RVT U58 ( .A1(n61), .A2(n24), .A3(n60), .A4(n21), .A5(n59), .A6(n43), 
        .Y(n74) );
  AO221X1_RVT U59 ( .A1(A[6]), .A2(n7), .A3(A[5]), .A4(n13), .A5(n75), .Y(n43)
         );
  AO22X1_RVT U60 ( .A1(A[7]), .A2(n11), .A3(A[8]), .A4(n10), .Y(n75) );
  AO221X1_RVT U61 ( .A1(A[10]), .A2(n7), .A3(A[9]), .A4(n13), .A5(n76), .Y(n21) );
  AO22X1_RVT U62 ( .A1(A[11]), .A2(n2), .A3(A[12]), .A4(n9), .Y(n76) );
  OA21X1_RVT U63 ( .A1(n77), .A2(n78), .A3(n54), .Y(n71) );
  AO22X1_RVT U64 ( .A1(A[1]), .A2(n13), .A3(A[2]), .A4(n8), .Y(n78) );
  AO22X1_RVT U65 ( .A1(A[3]), .A2(n2), .A3(A[4]), .A4(n9), .Y(n77) );
  AND3X1_RVT U66 ( .A1(n79), .A2(n63), .A3(n16), .Y(B[19]) );
  AND2X1_RVT U67 ( .A1(n66), .A2(n79), .Y(B[18]) );
  AND2X1_RVT U68 ( .A1(n16), .A2(n80), .Y(n66) );
  AND2X1_RVT U69 ( .A1(n73), .A2(n79), .Y(B[17]) );
  AND2X1_RVT U70 ( .A1(n16), .A2(n23), .Y(n73) );
  MUX21X1_RVT U71 ( .A1(n46), .A2(n45), .S0(n17), .Y(n23) );
  AND2X1_RVT U72 ( .A1(n81), .A2(n79), .Y(B[16]) );
  AO222X1_RVT U73 ( .A1(n20), .A2(n36), .A3(n35), .A4(n32), .A5(n1), .A6(n34), 
        .Y(B[15]) );
  AO222X1_RVT U74 ( .A1(n20), .A2(n40), .A3(n35), .A4(n42), .A5(n1), .A6(n41), 
        .Y(B[14]) );
  AO222X1_RVT U75 ( .A1(n20), .A2(n24), .A3(n35), .A4(n46), .A5(n1), .A6(n45), 
        .Y(B[13]) );
  AO221X1_RVT U76 ( .A1(A[18]), .A2(n8), .A3(A[17]), .A4(n13), .A5(n82), .Y(
        n45) );
  AO22X1_RVT U77 ( .A1(A[19]), .A2(n11), .A3(A[20]), .A4(n9), .Y(n82) );
  AO222X1_RVT U78 ( .A1(A[22]), .A2(n8), .A3(A[23]), .A4(n11), .A5(A[21]), 
        .A6(n12), .Y(n46) );
  AO221X1_RVT U79 ( .A1(A[14]), .A2(n7), .A3(A[13]), .A4(n13), .A5(n83), .Y(
        n24) );
  AO22X1_RVT U80 ( .A1(A[15]), .A2(n2), .A3(A[16]), .A4(n9), .Y(n83) );
  AO222X1_RVT U81 ( .A1(n20), .A2(n27), .A3(n35), .A4(n50), .A5(n1), .A6(n49), 
        .Y(B[12]) );
  AND2X1_RVT U82 ( .A1(n22), .A2(n17), .Y(n35) );
  AO222X1_RVT U83 ( .A1(n1), .A2(n36), .A3(n20), .A4(n29), .A5(n22), .A6(n63), 
        .Y(B[11]) );
  MUX21X1_RVT U84 ( .A1(n32), .A2(n34), .S0(n17), .Y(n63) );
  AO221X1_RVT U85 ( .A1(A[20]), .A2(n7), .A3(A[19]), .A4(n13), .A5(n84), .Y(
        n34) );
  AO22X1_RVT U86 ( .A1(A[21]), .A2(n11), .A3(n9), .A4(A[22]), .Y(n84) );
  AND2X1_RVT U87 ( .A1(n12), .A2(A[23]), .Y(n32) );
  AO221X1_RVT U88 ( .A1(A[12]), .A2(n7), .A3(A[11]), .A4(n12), .A5(n85), .Y(
        n29) );
  AO22X1_RVT U89 ( .A1(A[13]), .A2(n11), .A3(A[14]), .A4(n9), .Y(n85) );
  AO221X1_RVT U90 ( .A1(A[16]), .A2(n8), .A3(A[15]), .A4(n12), .A5(n86), .Y(
        n36) );
  AO22X1_RVT U91 ( .A1(A[17]), .A2(n11), .A3(A[18]), .A4(n10), .Y(n86) );
  AO222X1_RVT U92 ( .A1(n20), .A2(n38), .A3(n22), .A4(n80), .A5(n1), .A6(n40), 
        .Y(B[10]) );
  AO221X1_RVT U93 ( .A1(A[15]), .A2(n7), .A3(A[14]), .A4(n12), .A5(n87), .Y(
        n40) );
  AO22X1_RVT U94 ( .A1(A[16]), .A2(n11), .A3(A[17]), .A4(n9), .Y(n87) );
  MUX21X1_RVT U95 ( .A1(n42), .A2(n41), .S0(n17), .Y(n80) );
  AO221X1_RVT U96 ( .A1(A[19]), .A2(n8), .A3(A[18]), .A4(n12), .A5(n88), .Y(
        n41) );
  AO22X1_RVT U97 ( .A1(A[20]), .A2(n2), .A3(n10), .A4(A[21]), .Y(n88) );
  AO22X1_RVT U98 ( .A1(n13), .A2(A[22]), .A3(n8), .A4(A[23]), .Y(n42) );
  AND2X1_RVT U99 ( .A1(n79), .A2(n89), .Y(n22) );
  AND2X1_RVT U100 ( .A1(n15), .A2(n14), .Y(n79) );
  AO221X1_RVT U101 ( .A1(A[11]), .A2(n7), .A3(A[10]), .A4(n12), .A5(n90), .Y(
        n38) );
  AO22X1_RVT U102 ( .A1(A[12]), .A2(n11), .A3(A[13]), .A4(n9), .Y(n90) );
  OA21X1_RVT U103 ( .A1(n91), .A2(n92), .A3(n14), .Y(B[0]) );
  MUX21X1_RVT U104 ( .A1(n81), .A2(n93), .S0(n15), .Y(n92) );
  AO222X1_RVT U105 ( .A1(n61), .A2(n27), .A3(n60), .A4(n25), .A5(n59), .A6(n47), .Y(n93) );
  AO221X1_RVT U106 ( .A1(A[5]), .A2(n8), .A3(A[4]), .A4(n12), .A5(n94), .Y(n47) );
  AO22X1_RVT U107 ( .A1(A[6]), .A2(n11), .A3(A[7]), .A4(n10), .Y(n94) );
  AND2X1_RVT U108 ( .A1(n16), .A2(SH[2]), .Y(n59) );
  AO221X1_RVT U109 ( .A1(A[9]), .A2(n7), .A3(A[8]), .A4(n12), .A5(n95), .Y(n25) );
  AO22X1_RVT U110 ( .A1(A[10]), .A2(n2), .A3(A[11]), .A4(n9), .Y(n95) );
  AND2X1_RVT U111 ( .A1(n17), .A2(n89), .Y(n60) );
  AO221X1_RVT U112 ( .A1(A[13]), .A2(n8), .A3(A[12]), .A4(n12), .A5(n96), .Y(
        n27) );
  AO22X1_RVT U113 ( .A1(A[14]), .A2(n2), .A3(A[15]), .A4(n9), .Y(n96) );
  AND2X1_RVT U114 ( .A1(SH[2]), .A2(n89), .Y(n61) );
  AND2X1_RVT U115 ( .A1(n16), .A2(n26), .Y(n81) );
  MUX21X1_RVT U116 ( .A1(n50), .A2(n49), .S0(n17), .Y(n26) );
  AO221X1_RVT U117 ( .A1(A[17]), .A2(n8), .A3(A[16]), .A4(n12), .A5(n97), .Y(
        n49) );
  AO22X1_RVT U118 ( .A1(A[18]), .A2(n2), .A3(A[19]), .A4(n10), .Y(n97) );
  AO221X1_RVT U119 ( .A1(A[21]), .A2(n8), .A3(A[20]), .A4(n12), .A5(n98), .Y(
        n50) );
  AO22X1_RVT U120 ( .A1(A[22]), .A2(n11), .A3(n10), .A4(A[23]), .Y(n98) );
  OA21X1_RVT U121 ( .A1(n99), .A2(n100), .A3(n54), .Y(n91) );
  AND3X1_RVT U122 ( .A1(n15), .A2(n17), .A3(n16), .Y(n54) );
  OR2X1_RVT U123 ( .A1(SH[3]), .A2(n101), .Y(n89) );
  OR2X1_RVT U124 ( .A1(SH[4]), .A2(n101), .Y(n51) );
  OR2X1_RVT U125 ( .A1(SH[5]), .A2(SH[6]), .Y(n101) );
  AO22X1_RVT U126 ( .A1(A[0]), .A2(n13), .A3(A[1]), .A4(n8), .Y(n100) );
  AO22X1_RVT U127 ( .A1(A[2]), .A2(n2), .A3(A[3]), .A4(n9), .Y(n99) );
endmodule


module fpu_DW01_sub_28 ( A, B, CI, DIFF, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [9:0] carry;

  FADDX1_RVT U2_7 ( .A(A[7]), .B(n2), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n3), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1_RVT U2_4 ( .A(A[4]), .B(n5), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n4), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n6), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n7), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n8), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  INVX1_RVT U1 ( .A(B[1]), .Y(n8) );
  INVX1_RVT U2 ( .A(B[3]), .Y(n6) );
  INVX1_RVT U3 ( .A(B[2]), .Y(n7) );
  INVX1_RVT U4 ( .A(B[4]), .Y(n5) );
  INVX1_RVT U5 ( .A(B[5]), .Y(n4) );
  INVX1_RVT U6 ( .A(B[6]), .Y(n3) );
  INVX1_RVT U7 ( .A(B[7]), .Y(n2) );
  INVX1_RVT U8 ( .A(B[0]), .Y(n9) );
  INVX1_RVT U9 ( .A(carry[8]), .Y(DIFF[8]) );
  OR2X1_RVT U10 ( .A1(n9), .A2(A[0]), .Y(carry[1]) );
  XNOR2X1_RVT U11 ( .A1(A[0]), .A2(n9), .Y(DIFF[0]) );
endmodule


module fpu_DW01_add_5 ( A, B, CI, SUM, CO );
  input [24:0] A;
  input [24:0] B;
  output [24:0] SUM;
  input CI;
  output CO;

  wire   [24:1] carry;

  FADDX1_RVT U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(
        SUM[9]) );
  FADDX1_RVT U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1_RVT U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(
        SUM[8]) );
  FADDX1_RVT U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1_RVT U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1_RVT U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1_RVT U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1_RVT U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(
        SUM[6]) );
  FADDX1_RVT U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(
        SUM[7]) );
  FADDX1_RVT U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(
        SUM[5]) );
  FADDX1_RVT U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FADDX1_RVT U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(
        SUM[4]) );
  FADDX1_RVT U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(
        SUM[2]) );
  FADDX1_RVT U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(
        SUM[3]) );
  FADDX1_RVT U1_1 ( .A(A[1]), .B(B[1]), .CI(carry[1]), .CO(carry[2]), .S(
        SUM[1]) );
  FADDX1_RVT U1_22 ( .A(A[22]), .B(B[22]), .CI(carry[22]), .CO(carry[23]), .S(
        SUM[22]) );
  FADDX1_RVT U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .CO(carry[21]), .S(
        SUM[20]) );
  FADDX1_RVT U1_21 ( .A(A[21]), .B(B[21]), .CI(carry[21]), .CO(carry[22]), .S(
        SUM[21]) );
  FADDX1_RVT U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FADDX1_RVT U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FADDX1_RVT U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FADDX1_RVT U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FADDX1_RVT U1_23 ( .A(A[23]), .B(B[23]), .CI(carry[23]), .CO(SUM[24]), .S(
        SUM[23]) );
  AND2X1_RVT U1 ( .A1(A[0]), .A2(B[0]), .Y(carry[1]) );
  XOR2X1_RVT U2 ( .A1(A[0]), .A2(B[0]), .Y(SUM[0]) );
endmodule


module fpu_DW_rash_1 ( A, DATA_TC, SH, SH_TC, B );
  input [23:0] A;
  input [7:0] SH;
  output [23:0] B;
  input DATA_TC, SH_TC;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;

  INVX1_RVT U3 ( .A(SH[0]), .Y(n17) );
  AND2X1_RVT U4 ( .A1(n57), .A2(n77), .Y(n2) );
  AOI21X1_RVT U5 ( .A1(n50), .A2(n51), .A3(SH[7]), .Y(B[3]) );
  MUX21X1_RVT U6 ( .A1(n55), .A2(n56), .S0(n13), .Y(n50) );
  AND2X1_RVT U7 ( .A1(SH[0]), .A2(n16), .Y(n1) );
  INVX1_RVT U8 ( .A(n5), .Y(n6) );
  INVX1_RVT U9 ( .A(n7), .Y(n8) );
  INVX1_RVT U10 ( .A(n49), .Y(n13) );
  INVX1_RVT U11 ( .A(n87), .Y(n14) );
  INVX1_RVT U12 ( .A(n8), .Y(n9) );
  AND2X1_RVT U13 ( .A1(n17), .A2(SH[1]), .Y(n3) );
  INVX1_RVT U14 ( .A(n4), .Y(n11) );
  INVX1_RVT U15 ( .A(n4), .Y(n10) );
  NAND2X0_RVT U16 ( .A1(n17), .A2(n16), .Y(n4) );
  AND2X1_RVT U17 ( .A1(n52), .A2(n12), .Y(n18) );
  INVX1_RVT U18 ( .A(SH[1]), .Y(n16) );
  NAND2X0_RVT U19 ( .A1(SH[0]), .A2(n16), .Y(n5) );
  INVX1_RVT U20 ( .A(SH[2]), .Y(n15) );
  INVX1_RVT U21 ( .A(SH[7]), .Y(n12) );
  AND2X1_RVT U22 ( .A1(SH[0]), .A2(SH[1]), .Y(n7) );
  AO222X1_RVT U23 ( .A1(n18), .A2(n19), .A3(n20), .A4(n21), .A5(n2), .A6(n22), 
        .Y(B[9]) );
  AO222X1_RVT U24 ( .A1(n18), .A2(n23), .A3(n20), .A4(n24), .A5(n2), .A6(n25), 
        .Y(B[8]) );
  AO221X1_RVT U25 ( .A1(n18), .A2(n26), .A3(n2), .A4(n27), .A5(n28), .Y(B[7])
         );
  AO222X1_RVT U26 ( .A1(n29), .A2(n30), .A3(n31), .A4(n32), .A5(n33), .A6(n34), 
        .Y(n28) );
  AO221X1_RVT U27 ( .A1(n18), .A2(n35), .A3(n2), .A4(n36), .A5(n37), .Y(B[6])
         );
  AO222X1_RVT U28 ( .A1(n33), .A2(n38), .A3(n31), .A4(n39), .A5(n29), .A6(n40), 
        .Y(n37) );
  AO221X1_RVT U29 ( .A1(n18), .A2(n41), .A3(n2), .A4(n19), .A5(n42), .Y(B[5])
         );
  AO222X1_RVT U30 ( .A1(n33), .A2(n22), .A3(n31), .A4(n43), .A5(n29), .A6(n44), 
        .Y(n42) );
  AO221X1_RVT U31 ( .A1(n18), .A2(n45), .A3(n2), .A4(n23), .A5(n46), .Y(B[4])
         );
  AO222X1_RVT U32 ( .A1(n33), .A2(n25), .A3(n31), .A4(n47), .A5(n29), .A6(n48), 
        .Y(n46) );
  AND4X1_RVT U33 ( .A1(n14), .A2(n15), .A3(n49), .A4(n12), .Y(n29) );
  AND2X1_RVT U34 ( .A1(n20), .A2(SH[2]), .Y(n31) );
  NAND2X0_RVT U35 ( .A1(n52), .A2(n53), .Y(n51) );
  AO221X1_RVT U36 ( .A1(A[4]), .A2(n6), .A3(A[3]), .A4(n10), .A5(n54), .Y(n53)
         );
  AO22X1_RVT U37 ( .A1(A[5]), .A2(n3), .A3(A[6]), .A4(n7), .Y(n54) );
  AOI222X1_RVT U38 ( .A1(n26), .A2(n57), .A3(n27), .A4(n58), .A5(n34), .A6(n59), .Y(n56) );
  AO221X1_RVT U39 ( .A1(A[8]), .A2(n6), .A3(A[7]), .A4(n11), .A5(n60), .Y(n26)
         );
  AO22X1_RVT U40 ( .A1(A[9]), .A2(n3), .A3(A[10]), .A4(n7), .Y(n60) );
  NAND2X0_RVT U41 ( .A1(n14), .A2(n61), .Y(n55) );
  OA21X1_RVT U42 ( .A1(n62), .A2(n63), .A3(n12), .Y(B[2]) );
  MUX21X1_RVT U43 ( .A1(n64), .A2(n65), .S0(n13), .Y(n63) );
  AO222X1_RVT U44 ( .A1(n59), .A2(n38), .A3(n58), .A4(n36), .A5(n57), .A6(n35), 
        .Y(n65) );
  AO221X1_RVT U45 ( .A1(A[7]), .A2(n6), .A3(A[6]), .A4(n11), .A5(n66), .Y(n35)
         );
  AO22X1_RVT U46 ( .A1(A[8]), .A2(n3), .A3(A[9]), .A4(n9), .Y(n66) );
  OA21X1_RVT U47 ( .A1(n67), .A2(n68), .A3(n52), .Y(n62) );
  AO22X1_RVT U48 ( .A1(A[2]), .A2(n11), .A3(A[3]), .A4(n1), .Y(n68) );
  AO22X1_RVT U49 ( .A1(A[4]), .A2(n3), .A3(A[5]), .A4(n9), .Y(n67) );
  AND2X1_RVT U50 ( .A1(n30), .A2(n18), .Y(B[23]) );
  AND2X1_RVT U51 ( .A1(n18), .A2(n40), .Y(B[22]) );
  AND2X1_RVT U52 ( .A1(n18), .A2(n44), .Y(B[21]) );
  AND2X1_RVT U53 ( .A1(n18), .A2(n48), .Y(B[20]) );
  OA21X1_RVT U54 ( .A1(n69), .A2(n70), .A3(n12), .Y(B[1]) );
  MUX21X1_RVT U55 ( .A1(n71), .A2(n72), .S0(n13), .Y(n70) );
  AO222X1_RVT U56 ( .A1(n59), .A2(n22), .A3(n58), .A4(n19), .A5(n57), .A6(n41), 
        .Y(n72) );
  AO221X1_RVT U57 ( .A1(A[6]), .A2(n6), .A3(A[5]), .A4(n11), .A5(n73), .Y(n41)
         );
  AO22X1_RVT U58 ( .A1(A[7]), .A2(n3), .A3(A[8]), .A4(n9), .Y(n73) );
  AO221X1_RVT U59 ( .A1(A[10]), .A2(n6), .A3(A[9]), .A4(n11), .A5(n74), .Y(n19) );
  AO22X1_RVT U60 ( .A1(A[11]), .A2(n3), .A3(A[12]), .A4(n9), .Y(n74) );
  OA21X1_RVT U61 ( .A1(n75), .A2(n76), .A3(n52), .Y(n69) );
  AO22X1_RVT U62 ( .A1(A[1]), .A2(n11), .A3(A[2]), .A4(n1), .Y(n76) );
  AO22X1_RVT U63 ( .A1(A[3]), .A2(n3), .A3(A[4]), .A4(n9), .Y(n75) );
  AND3X1_RVT U64 ( .A1(n77), .A2(n61), .A3(n14), .Y(B[19]) );
  AND2X1_RVT U65 ( .A1(n64), .A2(n77), .Y(B[18]) );
  AND2X1_RVT U66 ( .A1(n14), .A2(n78), .Y(n64) );
  AND2X1_RVT U67 ( .A1(n71), .A2(n77), .Y(B[17]) );
  AND2X1_RVT U68 ( .A1(n14), .A2(n21), .Y(n71) );
  MUX21X1_RVT U69 ( .A1(n44), .A2(n43), .S0(n15), .Y(n21) );
  AND2X1_RVT U70 ( .A1(n79), .A2(n77), .Y(B[16]) );
  AO222X1_RVT U71 ( .A1(n18), .A2(n34), .A3(n33), .A4(n30), .A5(n2), .A6(n32), 
        .Y(B[15]) );
  AO222X1_RVT U72 ( .A1(n18), .A2(n38), .A3(n33), .A4(n40), .A5(n2), .A6(n39), 
        .Y(B[14]) );
  AO222X1_RVT U73 ( .A1(n18), .A2(n22), .A3(n33), .A4(n44), .A5(n2), .A6(n43), 
        .Y(B[13]) );
  AO221X1_RVT U74 ( .A1(A[18]), .A2(n6), .A3(A[17]), .A4(n11), .A5(n80), .Y(
        n43) );
  AO22X1_RVT U75 ( .A1(A[19]), .A2(n3), .A3(A[20]), .A4(n7), .Y(n80) );
  AO222X1_RVT U76 ( .A1(A[22]), .A2(n1), .A3(A[23]), .A4(n3), .A5(A[21]), .A6(
        n10), .Y(n44) );
  AO221X1_RVT U77 ( .A1(A[14]), .A2(n6), .A3(A[13]), .A4(n11), .A5(n81), .Y(
        n22) );
  AO22X1_RVT U78 ( .A1(A[15]), .A2(n3), .A3(A[16]), .A4(n9), .Y(n81) );
  AO222X1_RVT U79 ( .A1(n18), .A2(n25), .A3(n33), .A4(n48), .A5(n2), .A6(n47), 
        .Y(B[12]) );
  AND2X1_RVT U80 ( .A1(n20), .A2(n15), .Y(n33) );
  AO222X1_RVT U81 ( .A1(n2), .A2(n34), .A3(n18), .A4(n27), .A5(n20), .A6(n61), 
        .Y(B[11]) );
  MUX21X1_RVT U82 ( .A1(n30), .A2(n32), .S0(n15), .Y(n61) );
  AO221X1_RVT U83 ( .A1(A[20]), .A2(n6), .A3(A[19]), .A4(n11), .A5(n82), .Y(
        n32) );
  AO22X1_RVT U84 ( .A1(A[21]), .A2(n3), .A3(n9), .A4(A[22]), .Y(n82) );
  AND2X1_RVT U85 ( .A1(n10), .A2(A[23]), .Y(n30) );
  AO221X1_RVT U86 ( .A1(A[12]), .A2(n6), .A3(A[11]), .A4(n10), .A5(n83), .Y(
        n27) );
  AO22X1_RVT U87 ( .A1(A[13]), .A2(n3), .A3(A[14]), .A4(n9), .Y(n83) );
  AO221X1_RVT U88 ( .A1(A[16]), .A2(n6), .A3(A[15]), .A4(n10), .A5(n84), .Y(
        n34) );
  AO22X1_RVT U89 ( .A1(A[17]), .A2(n3), .A3(A[18]), .A4(n7), .Y(n84) );
  AO222X1_RVT U90 ( .A1(n18), .A2(n36), .A3(n20), .A4(n78), .A5(n2), .A6(n38), 
        .Y(B[10]) );
  AO221X1_RVT U91 ( .A1(A[15]), .A2(n6), .A3(A[14]), .A4(n10), .A5(n85), .Y(
        n38) );
  AO22X1_RVT U92 ( .A1(A[16]), .A2(n3), .A3(A[17]), .A4(n7), .Y(n85) );
  MUX21X1_RVT U93 ( .A1(n40), .A2(n39), .S0(n15), .Y(n78) );
  AO221X1_RVT U94 ( .A1(A[19]), .A2(n6), .A3(A[18]), .A4(n10), .A5(n86), .Y(
        n39) );
  AO22X1_RVT U95 ( .A1(A[20]), .A2(n3), .A3(n9), .A4(A[21]), .Y(n86) );
  AO22X1_RVT U96 ( .A1(n11), .A2(A[22]), .A3(n6), .A4(A[23]), .Y(n40) );
  AND2X1_RVT U97 ( .A1(n77), .A2(n87), .Y(n20) );
  AND2X1_RVT U98 ( .A1(n13), .A2(n12), .Y(n77) );
  AO221X1_RVT U99 ( .A1(A[11]), .A2(n6), .A3(A[10]), .A4(n10), .A5(n88), .Y(
        n36) );
  AO22X1_RVT U100 ( .A1(A[12]), .A2(n3), .A3(A[13]), .A4(n7), .Y(n88) );
  OA21X1_RVT U101 ( .A1(n89), .A2(n90), .A3(n12), .Y(B[0]) );
  MUX21X1_RVT U102 ( .A1(n79), .A2(n91), .S0(n13), .Y(n90) );
  AO222X1_RVT U103 ( .A1(n59), .A2(n25), .A3(n58), .A4(n23), .A5(n57), .A6(n45), .Y(n91) );
  AO221X1_RVT U104 ( .A1(A[5]), .A2(n1), .A3(A[4]), .A4(n10), .A5(n92), .Y(n45) );
  AO22X1_RVT U105 ( .A1(A[6]), .A2(n3), .A3(A[7]), .A4(n7), .Y(n92) );
  AND2X1_RVT U106 ( .A1(n14), .A2(SH[2]), .Y(n57) );
  AO221X1_RVT U107 ( .A1(A[9]), .A2(n1), .A3(A[8]), .A4(n10), .A5(n93), .Y(n23) );
  AO22X1_RVT U108 ( .A1(A[10]), .A2(n3), .A3(A[11]), .A4(n9), .Y(n93) );
  AND2X1_RVT U109 ( .A1(n15), .A2(n87), .Y(n58) );
  AO221X1_RVT U110 ( .A1(A[13]), .A2(n1), .A3(A[12]), .A4(n10), .A5(n94), .Y(
        n25) );
  AO22X1_RVT U111 ( .A1(A[14]), .A2(n3), .A3(A[15]), .A4(n7), .Y(n94) );
  AND2X1_RVT U112 ( .A1(SH[2]), .A2(n87), .Y(n59) );
  AND2X1_RVT U113 ( .A1(n14), .A2(n24), .Y(n79) );
  MUX21X1_RVT U114 ( .A1(n48), .A2(n47), .S0(n15), .Y(n24) );
  AO221X1_RVT U115 ( .A1(A[17]), .A2(n1), .A3(A[16]), .A4(n10), .A5(n95), .Y(
        n47) );
  AO22X1_RVT U116 ( .A1(A[18]), .A2(n3), .A3(A[19]), .A4(n7), .Y(n95) );
  AO221X1_RVT U117 ( .A1(A[21]), .A2(n1), .A3(A[20]), .A4(n10), .A5(n96), .Y(
        n48) );
  AO22X1_RVT U118 ( .A1(A[22]), .A2(n3), .A3(n7), .A4(A[23]), .Y(n96) );
  OA21X1_RVT U119 ( .A1(n97), .A2(n98), .A3(n52), .Y(n89) );
  AND3X1_RVT U120 ( .A1(n13), .A2(n15), .A3(n14), .Y(n52) );
  OR2X1_RVT U121 ( .A1(SH[3]), .A2(n99), .Y(n87) );
  OR2X1_RVT U122 ( .A1(SH[4]), .A2(n99), .Y(n49) );
  OR2X1_RVT U123 ( .A1(SH[5]), .A2(SH[6]), .Y(n99) );
  AO22X1_RVT U124 ( .A1(A[0]), .A2(n11), .A3(A[1]), .A4(n1), .Y(n98) );
  AO22X1_RVT U125 ( .A1(A[2]), .A2(n3), .A3(A[3]), .A4(n9), .Y(n97) );
endmodule


module fpu_DW01_sub_29 ( A, B, CI, DIFF, CO );
  input [7:0] A;
  input [7:0] B;
  output [7:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8;
  wire   [8:0] carry;

  FADDX1_RVT U2_7 ( .A(A[7]), .B(n1), .CI(carry[7]), .S(DIFF[7]) );
  FADDX1_RVT U2_5 ( .A(A[5]), .B(n3), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5]) );
  FADDX1_RVT U2_3 ( .A(A[3]), .B(n5), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3]) );
  FADDX1_RVT U2_6 ( .A(A[6]), .B(n2), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6]) );
  FADDX1_RVT U2_4 ( .A(A[4]), .B(n4), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4]) );
  FADDX1_RVT U2_2 ( .A(A[2]), .B(n6), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2]) );
  FADDX1_RVT U2_1 ( .A(A[1]), .B(n7), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1]) );
  FADDX1_RVT U2_0 ( .A(A[0]), .B(n8), .CI(1'b1), .CO(carry[1]), .S(DIFF[0]) );
  INVX0_RVT U1 ( .A(B[0]), .Y(n8) );
  INVX0_RVT U2 ( .A(B[1]), .Y(n7) );
  INVX0_RVT U3 ( .A(B[2]), .Y(n6) );
  INVX0_RVT U4 ( .A(B[4]), .Y(n4) );
  INVX0_RVT U5 ( .A(B[6]), .Y(n2) );
  INVX0_RVT U6 ( .A(B[3]), .Y(n5) );
  INVX0_RVT U7 ( .A(B[5]), .Y(n3) );
  INVX0_RVT U8 ( .A(B[7]), .Y(n1) );
endmodule


module fpu_DW01_add_6 ( A, B, CI, SUM, CO );
  input [45:0] A;
  input [45:0] B;
  output [45:0] SUM;
  input CI;
  output CO;
  wire   \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n2,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111;
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX1_RVT U2 ( .A(n105), .Y(n23) );
  INVX1_RVT U3 ( .A(n110), .Y(n25) );
  INVX1_RVT U4 ( .A(n95), .Y(n20) );
  INVX1_RVT U5 ( .A(n98), .Y(n21) );
  INVX1_RVT U6 ( .A(n108), .Y(n24) );
  INVX1_RVT U7 ( .A(n91), .Y(n19) );
  INVX1_RVT U8 ( .A(n31), .Y(n4) );
  INVX1_RVT U9 ( .A(n71), .Y(n14) );
  INVX1_RVT U10 ( .A(n67), .Y(n13) );
  INVX1_RVT U11 ( .A(n63), .Y(n12) );
  INVX1_RVT U12 ( .A(n59), .Y(n11) );
  INVX1_RVT U13 ( .A(n55), .Y(n10) );
  INVX1_RVT U14 ( .A(n51), .Y(n9) );
  INVX1_RVT U15 ( .A(n47), .Y(n8) );
  INVX1_RVT U16 ( .A(n43), .Y(n7) );
  INVX1_RVT U17 ( .A(n39), .Y(n6) );
  INVX1_RVT U18 ( .A(n35), .Y(n5) );
  INVX1_RVT U19 ( .A(n75), .Y(n15) );
  INVX1_RVT U20 ( .A(n79), .Y(n16) );
  INVX1_RVT U21 ( .A(n83), .Y(n17) );
  INVX1_RVT U22 ( .A(n87), .Y(n18) );
  INVX1_RVT U23 ( .A(n97), .Y(n22) );
  INVX1_RVT U24 ( .A(B[44]), .Y(n3) );
  INVX1_RVT U25 ( .A(A[44]), .Y(n2) );
  AND2X1_RVT U26 ( .A1(n111), .A2(n110), .Y(SUM[23]) );
  XNOR2X1_RVT U27 ( .A1(B[45]), .A2(n26), .Y(SUM[45]) );
  OA22X1_RVT U28 ( .A1(n27), .A2(n3), .A3(n28), .A4(n2), .Y(n26) );
  AND2X1_RVT U29 ( .A1(n28), .A2(n2), .Y(n27) );
  XNOR3X1_RVT U30 ( .A1(B[44]), .A2(A[44]), .A3(n28), .Y(SUM[44]) );
  OA21X1_RVT U31 ( .A1(n29), .A2(n4), .A3(n30), .Y(n28) );
  XOR2X1_RVT U32 ( .A1(n32), .A2(n29), .Y(SUM[43]) );
  OA21X1_RVT U33 ( .A1(n33), .A2(n5), .A3(n34), .Y(n29) );
  NAND2X0_RVT U34 ( .A1(n31), .A2(n30), .Y(n32) );
  NAND2X0_RVT U35 ( .A1(B[43]), .A2(A[43]), .Y(n30) );
  OR2X1_RVT U36 ( .A1(B[43]), .A2(A[43]), .Y(n31) );
  XOR2X1_RVT U37 ( .A1(n36), .A2(n33), .Y(SUM[42]) );
  OA21X1_RVT U38 ( .A1(n37), .A2(n6), .A3(n38), .Y(n33) );
  NAND2X0_RVT U39 ( .A1(n35), .A2(n34), .Y(n36) );
  NAND2X0_RVT U40 ( .A1(B[42]), .A2(A[42]), .Y(n34) );
  OR2X1_RVT U41 ( .A1(B[42]), .A2(A[42]), .Y(n35) );
  XOR2X1_RVT U42 ( .A1(n40), .A2(n37), .Y(SUM[41]) );
  OA21X1_RVT U43 ( .A1(n41), .A2(n7), .A3(n42), .Y(n37) );
  NAND2X0_RVT U44 ( .A1(n39), .A2(n38), .Y(n40) );
  NAND2X0_RVT U45 ( .A1(B[41]), .A2(A[41]), .Y(n38) );
  OR2X1_RVT U46 ( .A1(B[41]), .A2(A[41]), .Y(n39) );
  XOR2X1_RVT U47 ( .A1(n44), .A2(n41), .Y(SUM[40]) );
  OA21X1_RVT U48 ( .A1(n45), .A2(n8), .A3(n46), .Y(n41) );
  NAND2X0_RVT U49 ( .A1(n43), .A2(n42), .Y(n44) );
  NAND2X0_RVT U50 ( .A1(B[40]), .A2(A[40]), .Y(n42) );
  OR2X1_RVT U51 ( .A1(B[40]), .A2(A[40]), .Y(n43) );
  XOR2X1_RVT U52 ( .A1(n48), .A2(n45), .Y(SUM[39]) );
  OA21X1_RVT U53 ( .A1(n49), .A2(n9), .A3(n50), .Y(n45) );
  NAND2X0_RVT U54 ( .A1(n47), .A2(n46), .Y(n48) );
  NAND2X0_RVT U55 ( .A1(B[39]), .A2(A[39]), .Y(n46) );
  OR2X1_RVT U56 ( .A1(B[39]), .A2(A[39]), .Y(n47) );
  XOR2X1_RVT U57 ( .A1(n52), .A2(n49), .Y(SUM[38]) );
  OA21X1_RVT U58 ( .A1(n53), .A2(n10), .A3(n54), .Y(n49) );
  NAND2X0_RVT U59 ( .A1(n51), .A2(n50), .Y(n52) );
  NAND2X0_RVT U60 ( .A1(B[38]), .A2(A[38]), .Y(n50) );
  OR2X1_RVT U61 ( .A1(B[38]), .A2(A[38]), .Y(n51) );
  XOR2X1_RVT U62 ( .A1(n56), .A2(n53), .Y(SUM[37]) );
  OA21X1_RVT U63 ( .A1(n57), .A2(n11), .A3(n58), .Y(n53) );
  NAND2X0_RVT U64 ( .A1(n55), .A2(n54), .Y(n56) );
  NAND2X0_RVT U65 ( .A1(B[37]), .A2(A[37]), .Y(n54) );
  OR2X1_RVT U66 ( .A1(B[37]), .A2(A[37]), .Y(n55) );
  XOR2X1_RVT U67 ( .A1(n60), .A2(n57), .Y(SUM[36]) );
  OA21X1_RVT U68 ( .A1(n61), .A2(n12), .A3(n62), .Y(n57) );
  NAND2X0_RVT U69 ( .A1(n59), .A2(n58), .Y(n60) );
  NAND2X0_RVT U70 ( .A1(B[36]), .A2(A[36]), .Y(n58) );
  OR2X1_RVT U71 ( .A1(B[36]), .A2(A[36]), .Y(n59) );
  XOR2X1_RVT U72 ( .A1(n64), .A2(n61), .Y(SUM[35]) );
  OA21X1_RVT U73 ( .A1(n65), .A2(n13), .A3(n66), .Y(n61) );
  NAND2X0_RVT U74 ( .A1(n63), .A2(n62), .Y(n64) );
  NAND2X0_RVT U75 ( .A1(B[35]), .A2(A[35]), .Y(n62) );
  OR2X1_RVT U76 ( .A1(B[35]), .A2(A[35]), .Y(n63) );
  XOR2X1_RVT U77 ( .A1(n68), .A2(n65), .Y(SUM[34]) );
  OA21X1_RVT U78 ( .A1(n69), .A2(n14), .A3(n70), .Y(n65) );
  NAND2X0_RVT U79 ( .A1(n67), .A2(n66), .Y(n68) );
  NAND2X0_RVT U80 ( .A1(B[34]), .A2(A[34]), .Y(n66) );
  OR2X1_RVT U81 ( .A1(B[34]), .A2(A[34]), .Y(n67) );
  XOR2X1_RVT U82 ( .A1(n72), .A2(n69), .Y(SUM[33]) );
  OA21X1_RVT U83 ( .A1(n73), .A2(n15), .A3(n74), .Y(n69) );
  NAND2X0_RVT U84 ( .A1(n71), .A2(n70), .Y(n72) );
  NAND2X0_RVT U85 ( .A1(B[33]), .A2(A[33]), .Y(n70) );
  OR2X1_RVT U86 ( .A1(B[33]), .A2(A[33]), .Y(n71) );
  XOR2X1_RVT U87 ( .A1(n76), .A2(n73), .Y(SUM[32]) );
  OA21X1_RVT U88 ( .A1(n77), .A2(n16), .A3(n78), .Y(n73) );
  NAND2X0_RVT U89 ( .A1(n75), .A2(n74), .Y(n76) );
  NAND2X0_RVT U90 ( .A1(B[32]), .A2(A[32]), .Y(n74) );
  OR2X1_RVT U91 ( .A1(B[32]), .A2(A[32]), .Y(n75) );
  XOR2X1_RVT U92 ( .A1(n80), .A2(n77), .Y(SUM[31]) );
  OA21X1_RVT U93 ( .A1(n81), .A2(n17), .A3(n82), .Y(n77) );
  NAND2X0_RVT U94 ( .A1(n79), .A2(n78), .Y(n80) );
  NAND2X0_RVT U95 ( .A1(B[31]), .A2(A[31]), .Y(n78) );
  OR2X1_RVT U96 ( .A1(B[31]), .A2(A[31]), .Y(n79) );
  XOR2X1_RVT U97 ( .A1(n84), .A2(n81), .Y(SUM[30]) );
  OA21X1_RVT U98 ( .A1(n85), .A2(n18), .A3(n86), .Y(n81) );
  NAND2X0_RVT U99 ( .A1(n83), .A2(n82), .Y(n84) );
  NAND2X0_RVT U100 ( .A1(B[30]), .A2(A[30]), .Y(n82) );
  OR2X1_RVT U101 ( .A1(B[30]), .A2(A[30]), .Y(n83) );
  XOR2X1_RVT U102 ( .A1(n88), .A2(n85), .Y(SUM[29]) );
  AOI21X1_RVT U103 ( .A1(n89), .A2(n90), .A3(n19), .Y(n85) );
  NAND2X0_RVT U104 ( .A1(n87), .A2(n86), .Y(n88) );
  NAND2X0_RVT U105 ( .A1(B[29]), .A2(A[29]), .Y(n86) );
  OR2X1_RVT U106 ( .A1(B[29]), .A2(A[29]), .Y(n87) );
  XNOR2X1_RVT U107 ( .A1(n92), .A2(n89), .Y(SUM[28]) );
  AO21X1_RVT U108 ( .A1(n93), .A2(n94), .A3(n20), .Y(n89) );
  AO21X1_RVT U109 ( .A1(n96), .A2(n97), .A3(n21), .Y(n93) );
  AO21X1_RVT U110 ( .A1(n99), .A2(n100), .A3(n23), .Y(n96) );
  NAND2X0_RVT U111 ( .A1(n90), .A2(n91), .Y(n92) );
  NAND2X0_RVT U112 ( .A1(B[28]), .A2(A[28]), .Y(n91) );
  OR2X1_RVT U113 ( .A1(B[28]), .A2(A[28]), .Y(n90) );
  XOR2X1_RVT U114 ( .A1(n101), .A2(n102), .Y(SUM[27]) );
  OA21X1_RVT U115 ( .A1(n22), .A2(n103), .A3(n98), .Y(n102) );
  NAND2X0_RVT U116 ( .A1(n94), .A2(n95), .Y(n101) );
  NAND2X0_RVT U117 ( .A1(B[27]), .A2(A[27]), .Y(n95) );
  OR2X1_RVT U118 ( .A1(B[27]), .A2(A[27]), .Y(n94) );
  XOR2X1_RVT U119 ( .A1(n104), .A2(n103), .Y(SUM[26]) );
  AOI21X1_RVT U120 ( .A1(n99), .A2(n100), .A3(n23), .Y(n103) );
  NAND2X0_RVT U121 ( .A1(n97), .A2(n98), .Y(n104) );
  NAND2X0_RVT U122 ( .A1(B[26]), .A2(A[26]), .Y(n98) );
  OR2X1_RVT U123 ( .A1(B[26]), .A2(A[26]), .Y(n97) );
  XNOR2X1_RVT U124 ( .A1(n106), .A2(n99), .Y(SUM[25]) );
  AO21X1_RVT U125 ( .A1(n25), .A2(n107), .A3(n24), .Y(n99) );
  NAND2X0_RVT U126 ( .A1(n100), .A2(n105), .Y(n106) );
  NAND2X0_RVT U127 ( .A1(B[25]), .A2(A[25]), .Y(n105) );
  OR2X1_RVT U128 ( .A1(B[25]), .A2(A[25]), .Y(n100) );
  XNOR2X1_RVT U129 ( .A1(n109), .A2(n25), .Y(SUM[24]) );
  NAND2X0_RVT U130 ( .A1(n107), .A2(n108), .Y(n109) );
  NAND2X0_RVT U131 ( .A1(B[24]), .A2(A[24]), .Y(n108) );
  OR2X1_RVT U132 ( .A1(B[24]), .A2(A[24]), .Y(n107) );
  NAND2X0_RVT U133 ( .A1(B[23]), .A2(A[23]), .Y(n110) );
  OR2X1_RVT U134 ( .A1(B[23]), .A2(A[23]), .Y(n111) );
endmodule


module fpu_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [23:0] A;
  input [23:0] B;
  output [47:0] PRODUCT;
  input TC;
  wire   \ab[23][23] , \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] ,
         \ab[23][18] , \ab[23][17] , \ab[23][16] , \ab[23][15] , \ab[23][14] ,
         \ab[23][13] , \ab[23][12] , \ab[23][11] , \ab[23][10] , \ab[23][9] ,
         \ab[23][8] , \ab[23][7] , \ab[23][6] , \ab[23][5] , \ab[23][4] ,
         \ab[23][3] , \ab[23][2] , \ab[23][1] , \ab[23][0] , \ab[22][23] ,
         \ab[22][22] , \ab[22][21] , \ab[22][20] , \ab[22][19] , \ab[22][18] ,
         \ab[22][17] , \ab[22][16] , \ab[22][15] , \ab[22][14] , \ab[22][13] ,
         \ab[22][12] , \ab[22][11] , \ab[22][10] , \ab[22][9] , \ab[22][8] ,
         \ab[22][7] , \ab[22][6] , \ab[22][5] , \ab[22][4] , \ab[22][3] ,
         \ab[22][2] , \ab[22][1] , \ab[22][0] , \ab[21][23] , \ab[21][22] ,
         \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] ,
         \ab[21][16] , \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] ,
         \ab[21][11] , \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] ,
         \ab[21][6] , \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] ,
         \ab[21][1] , \ab[21][0] , \ab[20][23] , \ab[20][22] , \ab[20][21] ,
         \ab[20][20] , \ab[20][19] , \ab[20][18] , \ab[20][17] , \ab[20][16] ,
         \ab[20][15] , \ab[20][14] , \ab[20][13] , \ab[20][12] , \ab[20][11] ,
         \ab[20][10] , \ab[20][9] , \ab[20][8] , \ab[20][7] , \ab[20][6] ,
         \ab[20][5] , \ab[20][4] , \ab[20][3] , \ab[20][2] , \ab[20][1] ,
         \ab[20][0] , \ab[19][23] , \ab[19][22] , \ab[19][21] , \ab[19][20] ,
         \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] , \ab[19][15] ,
         \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] , \ab[19][10] ,
         \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] ,
         \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] ,
         \ab[18][23] , \ab[18][22] , \ab[18][21] , \ab[18][20] , \ab[18][19] ,
         \ab[18][18] , \ab[18][17] , \ab[18][16] , \ab[18][15] , \ab[18][14] ,
         \ab[18][13] , \ab[18][12] , \ab[18][11] , \ab[18][10] , \ab[18][9] ,
         \ab[18][8] , \ab[18][7] , \ab[18][6] , \ab[18][5] , \ab[18][4] ,
         \ab[18][3] , \ab[18][2] , \ab[18][1] , \ab[18][0] , \ab[17][23] ,
         \ab[17][22] , \ab[17][21] , \ab[17][20] , \ab[17][19] , \ab[17][18] ,
         \ab[17][17] , \ab[17][16] , \ab[17][15] , \ab[17][14] , \ab[17][13] ,
         \ab[17][12] , \ab[17][11] , \ab[17][10] , \ab[17][9] , \ab[17][8] ,
         \ab[17][7] , \ab[17][6] , \ab[17][5] , \ab[17][4] , \ab[17][3] ,
         \ab[17][2] , \ab[17][1] , \ab[17][0] , \ab[16][23] , \ab[16][22] ,
         \ab[16][21] , \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] ,
         \ab[16][16] , \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] ,
         \ab[16][11] , \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] ,
         \ab[16][6] , \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] ,
         \ab[16][1] , \ab[16][0] , \ab[15][23] , \ab[15][22] , \ab[15][21] ,
         \ab[15][20] , \ab[15][19] , \ab[15][18] , \ab[15][17] , \ab[15][16] ,
         \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][23] , \ab[14][22] , \ab[14][21] , \ab[14][20] ,
         \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] , \ab[14][15] ,
         \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] , \ab[14][10] ,
         \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] ,
         \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] ,
         \ab[13][23] , \ab[13][22] , \ab[13][21] , \ab[13][20] , \ab[13][19] ,
         \ab[13][18] , \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][14] ,
         \ab[13][13] , \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] ,
         \ab[13][8] , \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] ,
         \ab[13][3] , \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][23] ,
         \ab[12][22] , \ab[12][21] , \ab[12][20] , \ab[12][19] , \ab[12][18] ,
         \ab[12][17] , \ab[12][16] , \ab[12][15] , \ab[12][14] , \ab[12][13] ,
         \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] , \ab[12][8] ,
         \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] , \ab[12][3] ,
         \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][23] , \ab[11][22] ,
         \ab[11][21] , \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] ,
         \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] ,
         \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] ,
         \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] ,
         \ab[11][1] , \ab[11][0] , \ab[10][23] , \ab[10][22] , \ab[10][21] ,
         \ab[10][20] , \ab[10][19] , \ab[10][18] , \ab[10][17] , \ab[10][16] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][23] , \ab[9][22] , \ab[9][21] , \ab[9][20] ,
         \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] , \ab[9][15] ,
         \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] , \ab[9][10] ,
         \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] ,
         \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] ,
         \ab[8][23] , \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] ,
         \ab[8][18] , \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] ,
         \ab[8][13] , \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] ,
         \ab[8][8] , \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] ,
         \ab[8][3] , \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][23] ,
         \ab[7][22] , \ab[7][21] , \ab[7][20] , \ab[7][19] , \ab[7][18] ,
         \ab[7][17] , \ab[7][16] , \ab[7][15] , \ab[7][14] , \ab[7][13] ,
         \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] , \ab[7][8] ,
         \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] , \ab[7][3] ,
         \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][23] , \ab[6][22] ,
         \ab[6][21] , \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] ,
         \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] ,
         \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] ,
         \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] ,
         \ab[6][1] , \ab[6][0] , \ab[5][23] , \ab[5][22] , \ab[5][21] ,
         \ab[5][20] , \ab[5][19] , \ab[5][18] , \ab[5][17] , \ab[5][16] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][23] , \ab[4][22] , \ab[4][21] , \ab[4][20] ,
         \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] , \ab[4][15] ,
         \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] ,
         \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] ,
         \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] ,
         \ab[3][23] , \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] ,
         \ab[3][18] , \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] ,
         \ab[3][13] , \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] ,
         \ab[3][8] , \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] ,
         \ab[3][3] , \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][23] ,
         \ab[2][22] , \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] ,
         \ab[2][17] , \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] ,
         \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][23] , \ab[1][22] ,
         \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] ,
         \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[1][0] , \ab[0][23] , \ab[0][22] , \ab[0][21] ,
         \ab[0][20] , \ab[0][19] , \ab[0][18] , \ab[0][17] , \ab[0][16] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[23][22] , \CARRYB[23][21] , \CARRYB[23][20] ,
         \CARRYB[23][19] , \CARRYB[23][18] , \CARRYB[23][17] ,
         \CARRYB[23][16] , \CARRYB[23][15] , \CARRYB[23][14] ,
         \CARRYB[23][13] , \CARRYB[23][12] , \CARRYB[23][11] ,
         \CARRYB[23][10] , \CARRYB[23][9] , \CARRYB[23][8] , \CARRYB[23][7] ,
         \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] , \CARRYB[23][3] ,
         \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][12] , \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] ,
         \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][22] , \CARRYB[21][21] , \CARRYB[21][20] ,
         \CARRYB[21][19] , \CARRYB[21][18] , \CARRYB[21][17] ,
         \CARRYB[21][16] , \CARRYB[21][15] , \CARRYB[21][14] ,
         \CARRYB[21][13] , \CARRYB[21][12] , \CARRYB[21][11] ,
         \CARRYB[21][10] , \CARRYB[21][9] , \CARRYB[21][8] , \CARRYB[21][7] ,
         \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] , \CARRYB[21][3] ,
         \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][22] , \CARRYB[19][21] , \CARRYB[19][20] ,
         \CARRYB[19][19] , \CARRYB[19][18] , \CARRYB[19][17] ,
         \CARRYB[19][16] , \CARRYB[19][15] , \CARRYB[19][14] ,
         \CARRYB[19][13] , \CARRYB[19][12] , \CARRYB[19][11] ,
         \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] , \CARRYB[19][7] ,
         \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] , \CARRYB[19][3] ,
         \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][22] , \CARRYB[17][21] , \CARRYB[17][20] ,
         \CARRYB[17][19] , \CARRYB[17][18] , \CARRYB[17][17] ,
         \CARRYB[17][16] , \CARRYB[17][15] , \CARRYB[17][14] ,
         \CARRYB[17][13] , \CARRYB[17][12] , \CARRYB[17][11] ,
         \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] , \CARRYB[17][7] ,
         \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] , \CARRYB[17][3] ,
         \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \CARRYB[15][22] , \CARRYB[15][21] , \CARRYB[15][20] ,
         \CARRYB[15][19] , \CARRYB[15][18] , \CARRYB[15][17] ,
         \CARRYB[15][16] , \CARRYB[15][15] , \CARRYB[15][14] ,
         \CARRYB[15][13] , \CARRYB[15][12] , \CARRYB[15][11] ,
         \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] , \CARRYB[15][7] ,
         \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][22] , \CARRYB[13][21] , \CARRYB[13][20] ,
         \CARRYB[13][19] , \CARRYB[13][18] , \CARRYB[13][17] ,
         \CARRYB[13][16] , \CARRYB[13][15] , \CARRYB[13][14] ,
         \CARRYB[13][13] , \CARRYB[13][12] , \CARRYB[13][11] ,
         \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] , \CARRYB[13][7] ,
         \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] , \CARRYB[13][3] ,
         \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][22] , \CARRYB[11][21] , \CARRYB[11][20] ,
         \CARRYB[11][19] , \CARRYB[11][18] , \CARRYB[11][17] ,
         \CARRYB[11][16] , \CARRYB[11][15] , \CARRYB[11][14] ,
         \CARRYB[11][13] , \CARRYB[11][12] , \CARRYB[11][11] ,
         \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] , \CARRYB[11][7] ,
         \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] , \CARRYB[11][3] ,
         \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] , \CARRYB[10][22] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][22] , \CARRYB[9][21] , \CARRYB[9][20] ,
         \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] , \CARRYB[9][16] ,
         \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] ,
         \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] ,
         \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] ,
         \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] ,
         \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] , \CARRYB[8][19] ,
         \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] ,
         \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] ,
         \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] ,
         \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][22] ,
         \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] ,
         \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][22] , \CARRYB[5][21] , \CARRYB[5][20] ,
         \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] , \CARRYB[5][16] ,
         \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] ,
         \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] ,
         \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] ,
         \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] ,
         \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] ,
         \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] ,
         \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] ,
         \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] ,
         \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] ,
         \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][22] , \CARRYB[2][21] ,
         \CARRYB[2][20] , \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] ,
         \CARRYB[2][16] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][22] , \CARRYB[1][21] , \CARRYB[1][20] ,
         \CARRYB[1][19] , \CARRYB[1][18] , \CARRYB[1][17] , \CARRYB[1][16] ,
         \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] , \CARRYB[1][12] ,
         \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][8] ,
         \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] ,
         \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] ,
         \SUMB[23][22] , \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] ,
         \SUMB[23][18] , \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] ,
         \SUMB[23][14] , \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] ,
         \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] ,
         \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] ,
         \SUMB[23][2] , \SUMB[23][1] , \SUMB[23][0] , \SUMB[22][22] ,
         \SUMB[22][21] , \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] ,
         \SUMB[22][17] , \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] ,
         \SUMB[22][13] , \SUMB[22][12] , \SUMB[22][11] , \SUMB[22][10] ,
         \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] , \SUMB[22][6] ,
         \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] , \SUMB[22][2] ,
         \SUMB[22][1] , \SUMB[21][22] , \SUMB[21][21] , \SUMB[21][20] ,
         \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] , \SUMB[21][16] ,
         \SUMB[21][15] , \SUMB[21][14] , \SUMB[21][13] , \SUMB[21][12] ,
         \SUMB[21][11] , \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] ,
         \SUMB[21][7] , \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] ,
         \SUMB[21][3] , \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][22] ,
         \SUMB[20][21] , \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] ,
         \SUMB[20][17] , \SUMB[20][16] , \SUMB[20][15] , \SUMB[20][14] ,
         \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] , \SUMB[20][10] ,
         \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] , \SUMB[20][6] ,
         \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] , \SUMB[20][2] ,
         \SUMB[20][1] , \SUMB[19][22] , \SUMB[19][21] , \SUMB[19][20] ,
         \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] , \SUMB[19][16] ,
         \SUMB[19][15] , \SUMB[19][14] , \SUMB[19][13] , \SUMB[19][12] ,
         \SUMB[19][11] , \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] ,
         \SUMB[19][7] , \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] ,
         \SUMB[19][3] , \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][22] ,
         \SUMB[18][21] , \SUMB[18][20] , \SUMB[18][19] , \SUMB[18][18] ,
         \SUMB[18][17] , \SUMB[18][16] , \SUMB[18][15] , \SUMB[18][14] ,
         \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] , \SUMB[18][10] ,
         \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] ,
         \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] ,
         \SUMB[18][1] , \SUMB[17][22] , \SUMB[17][21] , \SUMB[17][20] ,
         \SUMB[17][19] , \SUMB[17][18] , \SUMB[17][17] , \SUMB[17][16] ,
         \SUMB[17][15] , \SUMB[17][14] , \SUMB[17][13] , \SUMB[17][12] ,
         \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] , \SUMB[17][8] ,
         \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] ,
         \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][22] ,
         \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][19] , \SUMB[16][18] ,
         \SUMB[16][17] , \SUMB[16][16] , \SUMB[16][15] , \SUMB[16][14] ,
         \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][10] ,
         \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] ,
         \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] ,
         \SUMB[16][1] , \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] ,
         \SUMB[15][19] , \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] ,
         \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] ,
         \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] ,
         \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] ,
         \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][22] ,
         \SUMB[14][21] , \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] ,
         \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] ,
         \SUMB[13][19] , \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] ,
         \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][22] ,
         \SUMB[12][21] , \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] ,
         \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] ,
         \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] ,
         \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][22] ,
         \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] ,
         \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] ,
         \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] ,
         \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][22] , \SUMB[8][21] ,
         \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] , \SUMB[8][17] ,
         \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][22] ,
         \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] , \SUMB[6][18] ,
         \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][22] ,
         \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] , \SUMB[5][18] ,
         \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][22] ,
         \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] , \SUMB[4][18] ,
         \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][22] ,
         \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] ,
         \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[44] ,
         \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] ,
         \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] ,
         \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] ,
         \A1[22] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] ,
         \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] ,
         \A2[32] , \A2[31] , \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] ,
         \A2[25] , \A2[24] , \A2[23] , n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146;

  fpu_DW01_add_6 FS_1 ( .A({1'b0, \A1[44] , \A1[43] , \A1[42] , \A1[41] , 
        \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , 
        \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \SUMB[23][0] , 
        \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , 
        \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , 
        \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({
        \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , 
        \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , 
        \A2[31] , \A2[30] , \A2[29] , \A2[28] , \A2[27] , \A2[26] , \A2[25] , 
        \A2[24] , \A2[23] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[47:2]) );
  FADDX1_RVT S3_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(
        \ab[21][23] ), .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FADDX1_RVT S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(
        \SUMB[21][22] ), .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FADDX1_RVT S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(
        \SUMB[21][21] ), .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FADDX1_RVT S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(
        \SUMB[21][20] ), .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FADDX1_RVT S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(
        \SUMB[21][19] ), .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FADDX1_RVT S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(
        \SUMB[21][18] ), .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FADDX1_RVT S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(
        \SUMB[21][17] ), .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FADDX1_RVT S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(
        \SUMB[21][16] ), .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FADDX1_RVT S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(
        \SUMB[21][15] ), .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FADDX1_RVT S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(
        \SUMB[21][14] ), .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FADDX1_RVT S3_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(
        \ab[13][23] ), .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FADDX1_RVT S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(
        \SUMB[13][22] ), .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FADDX1_RVT S3_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(
        \ab[14][23] ), .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FADDX1_RVT S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(
        \SUMB[14][22] ), .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FADDX1_RVT S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(
        \SUMB[14][21] ), .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FADDX1_RVT S3_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(
        \ab[12][23] ), .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FADDX1_RVT S3_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(
        \ab[19][23] ), .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FADDX1_RVT S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(
        \SUMB[19][22] ), .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FADDX1_RVT S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(
        \SUMB[19][21] ), .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FADDX1_RVT S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(
        \SUMB[19][20] ), .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FADDX1_RVT S3_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(
        \ab[17][23] ), .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FADDX1_RVT S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(
        \SUMB[19][19] ), .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FADDX1_RVT S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(
        \SUMB[17][22] ), .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FADDX1_RVT S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(
        \SUMB[19][18] ), .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FADDX1_RVT S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(
        \SUMB[17][21] ), .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FADDX1_RVT S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(
        \SUMB[19][17] ), .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FADDX1_RVT S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(
        \SUMB[17][20] ), .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FADDX1_RVT S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(
        \SUMB[19][16] ), .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FADDX1_RVT S3_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(
        \ab[15][23] ), .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FADDX1_RVT S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(
        \SUMB[17][19] ), .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FADDX1_RVT S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(
        \SUMB[15][22] ), .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FADDX1_RVT S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(
        \SUMB[17][18] ), .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FADDX1_RVT S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(
        \SUMB[15][21] ), .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FADDX1_RVT S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(
        \SUMB[15][20] ), .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FADDX1_RVT S3_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(
        \ab[18][23] ), .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FADDX1_RVT S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(
        \SUMB[18][22] ), .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FADDX1_RVT S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(
        \SUMB[18][21] ), .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FADDX1_RVT S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(
        \SUMB[18][20] ), .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FADDX1_RVT S3_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(
        \ab[16][23] ), .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FADDX1_RVT S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(
        \SUMB[18][19] ), .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FADDX1_RVT S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(
        \SUMB[16][22] ), .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FADDX1_RVT S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(
        \SUMB[18][18] ), .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FADDX1_RVT S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(
        \SUMB[16][21] ), .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FADDX1_RVT S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(
        \SUMB[18][17] ), .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FADDX1_RVT S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(
        \SUMB[16][20] ), .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FADDX1_RVT S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(
        \SUMB[16][19] ), .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FADDX1_RVT S3_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(
        \ab[20][23] ), .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FADDX1_RVT S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(
        \SUMB[20][22] ), .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FADDX1_RVT S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(
        \SUMB[20][21] ), .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FADDX1_RVT S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(
        \SUMB[20][20] ), .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FADDX1_RVT S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(
        \SUMB[20][19] ), .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FADDX1_RVT S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(
        \SUMB[20][18] ), .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FADDX1_RVT S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(
        \SUMB[20][17] ), .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FADDX1_RVT S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(
        \SUMB[20][16] ), .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FADDX1_RVT S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(
        \SUMB[20][15] ), .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FADDX1_RVT S5_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\ab[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FADDX1_RVT S4_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(
        \SUMB[22][22] ), .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FADDX1_RVT S4_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(
        \SUMB[22][21] ), .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FADDX1_RVT S4_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(
        \SUMB[22][20] ), .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FADDX1_RVT S4_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(
        \SUMB[22][19] ), .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FADDX1_RVT S4_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(
        \SUMB[22][18] ), .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FADDX1_RVT S4_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(
        \SUMB[22][17] ), .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FADDX1_RVT S4_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(
        \SUMB[22][16] ), .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FADDX1_RVT S4_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(
        \SUMB[22][15] ), .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FADDX1_RVT S4_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(
        \SUMB[22][14] ), .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FADDX1_RVT S4_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(
        \SUMB[22][13] ), .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FADDX1_RVT S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FADDX1_RVT S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FADDX1_RVT S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FADDX1_RVT S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FADDX1_RVT S3_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\ab[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FADDX1_RVT S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FADDX1_RVT S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FADDX1_RVT S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(
        \SUMB[21][13] ), .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FADDX1_RVT S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(
        \SUMB[21][12] ), .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FADDX1_RVT S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(
        \SUMB[21][11] ), .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FADDX1_RVT S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(
        \SUMB[21][10] ), .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FADDX1_RVT S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FADDX1_RVT S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FADDX1_RVT S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FADDX1_RVT S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FADDX1_RVT S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FADDX1_RVT S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FADDX1_RVT S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FADDX1_RVT S3_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\ab[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FADDX1_RVT S3_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\ab[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FADDX1_RVT S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FADDX1_RVT S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FADDX1_RVT S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FADDX1_RVT S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FADDX1_RVT S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FADDX1_RVT S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FADDX1_RVT S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FADDX1_RVT S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FADDX1_RVT S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FADDX1_RVT S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FADDX1_RVT S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FADDX1_RVT S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FADDX1_RVT S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FADDX1_RVT S3_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\ab[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FADDX1_RVT S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FADDX1_RVT S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FADDX1_RVT S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FADDX1_RVT S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FADDX1_RVT S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FADDX1_RVT S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FADDX1_RVT S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(
        \SUMB[13][21] ), .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FADDX1_RVT S2_14_19 ( .A(\ab[14][19] ), .B(\CARRYB[13][19] ), .CI(
        \SUMB[13][20] ), .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FADDX1_RVT S3_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(
        \ab[11][23] ), .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FADDX1_RVT S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(
        \SUMB[13][19] ), .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FADDX1_RVT S2_12_21 ( .A(\ab[12][21] ), .B(\CARRYB[11][21] ), .CI(
        \SUMB[11][22] ), .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FADDX1_RVT S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(
        \SUMB[13][18] ), .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FADDX1_RVT S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(
        \SUMB[11][21] ), .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FADDX1_RVT S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(
        \SUMB[13][17] ), .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FADDX1_RVT S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(
        \SUMB[11][20] ), .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FADDX1_RVT S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(
        \SUMB[13][13] ), .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FADDX1_RVT S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(
        \SUMB[13][14] ), .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FADDX1_RVT S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(
        \SUMB[13][15] ), .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FADDX1_RVT S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(
        \SUMB[13][16] ), .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FADDX1_RVT S3_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\ab[9][23] ), .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FADDX1_RVT S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(
        \SUMB[11][19] ), .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FADDX1_RVT S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(
        \SUMB[9][22] ), .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FADDX1_RVT S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(
        \SUMB[11][15] ), .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FADDX1_RVT S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(
        \SUMB[11][16] ), .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FADDX1_RVT S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(
        \SUMB[11][17] ), .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FADDX1_RVT S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(
        \SUMB[11][18] ), .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FADDX1_RVT S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(
        \SUMB[9][21] ), .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FADDX1_RVT S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FADDX1_RVT S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FADDX1_RVT S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FADDX1_RVT S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(
        \SUMB[13][10] ), .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FADDX1_RVT S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(
        \SUMB[13][11] ), .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FADDX1_RVT S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(
        \SUMB[13][12] ), .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FADDX1_RVT S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(
        \SUMB[9][17] ), .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FADDX1_RVT S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(
        \SUMB[9][18] ), .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FADDX1_RVT S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(
        \SUMB[9][19] ), .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FADDX1_RVT S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(
        \SUMB[9][20] ), .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FADDX1_RVT S3_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\ab[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FADDX1_RVT S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FADDX1_RVT S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(
        \SUMB[11][10] ), .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FADDX1_RVT S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(
        \SUMB[11][11] ), .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FADDX1_RVT S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(
        \SUMB[11][12] ), .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FADDX1_RVT S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(
        \SUMB[11][13] ), .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FADDX1_RVT S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(
        \SUMB[11][14] ), .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FADDX1_RVT S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FADDX1_RVT S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FADDX1_RVT S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FADDX1_RVT S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FADDX1_RVT S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(
        \SUMB[9][11] ), .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FADDX1_RVT S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(
        \SUMB[9][12] ), .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FADDX1_RVT S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(
        \SUMB[9][13] ), .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FADDX1_RVT S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(
        \SUMB[9][14] ), .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FADDX1_RVT S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(
        \SUMB[9][15] ), .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FADDX1_RVT S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(
        \SUMB[9][16] ), .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FADDX1_RVT S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FADDX1_RVT S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FADDX1_RVT S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FADDX1_RVT S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FADDX1_RVT S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FADDX1_RVT S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FADDX1_RVT S2_15_19 ( .A(\ab[15][19] ), .B(\CARRYB[14][19] ), .CI(
        \SUMB[14][20] ), .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FADDX1_RVT S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(
        \SUMB[14][19] ), .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FADDX1_RVT S2_13_21 ( .A(\ab[13][21] ), .B(\CARRYB[12][21] ), .CI(
        \SUMB[12][22] ), .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FADDX1_RVT S2_15_17 ( .A(\ab[15][17] ), .B(\CARRYB[14][17] ), .CI(
        \SUMB[14][18] ), .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FADDX1_RVT S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(
        \SUMB[12][21] ), .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FADDX1_RVT S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(
        \SUMB[14][17] ), .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FADDX1_RVT S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(
        \SUMB[12][20] ), .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FADDX1_RVT S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(
        \SUMB[14][16] ), .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FADDX1_RVT S3_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(
        \ab[10][23] ), .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FADDX1_RVT S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(
        \SUMB[12][19] ), .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FADDX1_RVT S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(
        \SUMB[14][12] ), .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FADDX1_RVT S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(
        \SUMB[14][13] ), .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FADDX1_RVT S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(
        \SUMB[14][14] ), .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FADDX1_RVT S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(
        \SUMB[14][15] ), .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FADDX1_RVT S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(
        \SUMB[10][22] ), .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FADDX1_RVT S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(
        \SUMB[12][18] ), .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FADDX1_RVT S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(
        \SUMB[10][21] ), .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FADDX1_RVT S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(
        \SUMB[12][14] ), .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FADDX1_RVT S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(
        \SUMB[12][15] ), .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FADDX1_RVT S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(
        \SUMB[12][16] ), .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FADDX1_RVT S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(
        \SUMB[12][17] ), .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FADDX1_RVT S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(
        \SUMB[10][20] ), .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FADDX1_RVT S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FADDX1_RVT S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FADDX1_RVT S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FADDX1_RVT S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FADDX1_RVT S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(
        \SUMB[14][10] ), .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FADDX1_RVT S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(
        \SUMB[14][11] ), .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FADDX1_RVT S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(
        \SUMB[10][16] ), .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FADDX1_RVT S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(
        \SUMB[10][17] ), .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FADDX1_RVT S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(
        \SUMB[10][18] ), .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FADDX1_RVT S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(
        \SUMB[10][19] ), .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FADDX1_RVT S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FADDX1_RVT S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FADDX1_RVT S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(
        \SUMB[12][10] ), .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FADDX1_RVT S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(
        \SUMB[12][11] ), .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FADDX1_RVT S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(
        \SUMB[12][12] ), .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FADDX1_RVT S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(
        \SUMB[12][13] ), .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FADDX1_RVT S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(
        \SUMB[10][10] ), .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FADDX1_RVT S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(
        \SUMB[10][11] ), .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FADDX1_RVT S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(
        \SUMB[10][12] ), .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FADDX1_RVT S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(
        \SUMB[10][13] ), .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FADDX1_RVT S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(
        \SUMB[10][14] ), .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FADDX1_RVT S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(
        \SUMB[10][15] ), .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FADDX1_RVT S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FADDX1_RVT S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FADDX1_RVT S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FADDX1_RVT S3_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\ab[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FADDX1_RVT S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FADDX1_RVT S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FADDX1_RVT S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FADDX1_RVT S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FADDX1_RVT S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FADDX1_RVT S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FADDX1_RVT S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FADDX1_RVT S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(
        \SUMB[19][15] ), .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FADDX1_RVT S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(
        \SUMB[19][14] ), .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FADDX1_RVT S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(
        \SUMB[17][17] ), .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FADDX1_RVT S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(
        \SUMB[19][13] ), .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FADDX1_RVT S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(
        \SUMB[17][16] ), .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FADDX1_RVT S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(
        \SUMB[19][12] ), .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FADDX1_RVT S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(
        \SUMB[15][19] ), .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FADDX1_RVT S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(
        \SUMB[17][15] ), .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FADDX1_RVT S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(
        \SUMB[19][11] ), .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FADDX1_RVT S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(
        \SUMB[15][18] ), .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FADDX1_RVT S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(
        \SUMB[17][14] ), .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FADDX1_RVT S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FADDX1_RVT S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FADDX1_RVT S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(
        \SUMB[19][10] ), .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FADDX1_RVT S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FADDX1_RVT S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(
        \SUMB[15][17] ), .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FADDX1_RVT S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(
        \SUMB[17][13] ), .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FADDX1_RVT S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(
        \SUMB[15][16] ), .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FADDX1_RVT S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FADDX1_RVT S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(
        \SUMB[17][10] ), .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FADDX1_RVT S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(
        \SUMB[17][11] ), .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FADDX1_RVT S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(
        \SUMB[17][12] ), .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FADDX1_RVT S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(
        \SUMB[15][15] ), .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FADDX1_RVT S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FADDX1_RVT S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FADDX1_RVT S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FADDX1_RVT S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(
        \SUMB[15][11] ), .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FADDX1_RVT S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(
        \SUMB[15][12] ), .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FADDX1_RVT S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(
        \SUMB[15][13] ), .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FADDX1_RVT S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(
        \SUMB[15][14] ), .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FADDX1_RVT S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FADDX1_RVT S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FADDX1_RVT S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FADDX1_RVT S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FADDX1_RVT S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FADDX1_RVT S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FADDX1_RVT S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FADDX1_RVT S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FADDX1_RVT S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FADDX1_RVT S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FADDX1_RVT S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(
        \SUMB[15][10] ), .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FADDX1_RVT S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FADDX1_RVT S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(
        \SUMB[18][16] ), .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FADDX1_RVT S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(
        \SUMB[18][15] ), .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FADDX1_RVT S2_17_17 ( .A(\ab[17][17] ), .B(\CARRYB[16][17] ), .CI(
        \SUMB[16][18] ), .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FADDX1_RVT S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(
        \SUMB[18][14] ), .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FADDX1_RVT S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(
        \SUMB[16][17] ), .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FADDX1_RVT S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(
        \SUMB[18][13] ), .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FADDX1_RVT S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(
        \SUMB[16][16] ), .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FADDX1_RVT S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(
        \SUMB[18][12] ), .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FADDX1_RVT S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(
        \SUMB[16][15] ), .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FADDX1_RVT S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FADDX1_RVT S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FADDX1_RVT S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(
        \SUMB[18][10] ), .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FADDX1_RVT S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(
        \SUMB[18][11] ), .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FADDX1_RVT S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(
        \SUMB[16][14] ), .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FADDX1_RVT S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(
        \SUMB[16][10] ), .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FADDX1_RVT S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(
        \SUMB[16][11] ), .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FADDX1_RVT S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(
        \SUMB[16][12] ), .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FADDX1_RVT S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(
        \SUMB[16][13] ), .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FADDX1_RVT S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FADDX1_RVT S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FADDX1_RVT S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FADDX1_RVT S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FADDX1_RVT S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FADDX1_RVT S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FADDX1_RVT S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FADDX1_RVT S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FADDX1_RVT S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FADDX1_RVT S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FADDX1_RVT S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FADDX1_RVT S2_21_13 ( .A(\ab[21][13] ), .B(\CARRYB[20][13] ), .CI(
        \SUMB[20][14] ), .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FADDX1_RVT S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(
        \SUMB[20][13] ), .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FADDX1_RVT S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(
        \SUMB[20][12] ), .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FADDX1_RVT S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(
        \SUMB[20][11] ), .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FADDX1_RVT S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(
        \SUMB[20][10] ), .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FADDX1_RVT S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FADDX1_RVT S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FADDX1_RVT S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FADDX1_RVT S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FADDX1_RVT S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FADDX1_RVT S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FADDX1_RVT S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FADDX1_RVT S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FADDX1_RVT S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FADDX1_RVT S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FADDX1_RVT S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FADDX1_RVT S3_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\ab[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FADDX1_RVT S3_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\ab[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FADDX1_RVT S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FADDX1_RVT S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FADDX1_RVT S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FADDX1_RVT S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FADDX1_RVT S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FADDX1_RVT S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FADDX1_RVT S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FADDX1_RVT S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FADDX1_RVT S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FADDX1_RVT S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FADDX1_RVT S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FADDX1_RVT S4_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FADDX1_RVT S4_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FADDX1_RVT S4_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FADDX1_RVT S4_11 ( .A(\ab[23][11] ), .B(\CARRYB[22][11] ), .CI(
        \SUMB[22][12] ), .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FADDX1_RVT S4_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(
        \SUMB[22][11] ), .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FADDX1_RVT S4_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FADDX1_RVT S4_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FADDX1_RVT S4_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FADDX1_RVT S4_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FADDX1_RVT S4_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FADDX1_RVT S4_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\SUMB[23][0] ) );
  FADDX1_RVT S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FADDX1_RVT S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FADDX1_RVT S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FADDX1_RVT S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FADDX1_RVT S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FADDX1_RVT S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FADDX1_RVT S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FADDX1_RVT S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FADDX1_RVT S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FADDX1_RVT S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FADDX1_RVT S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FADDX1_RVT S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FADDX1_RVT S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FADDX1_RVT S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FADDX1_RVT S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FADDX1_RVT S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FADDX1_RVT S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FADDX1_RVT S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FADDX1_RVT S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FADDX1_RVT S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FADDX1_RVT S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FADDX1_RVT S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FADDX1_RVT S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), 
        .CO(\CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FADDX1_RVT S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), 
        .CO(\CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FADDX1_RVT S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FADDX1_RVT S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FADDX1_RVT S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), 
        .CO(\CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FADDX1_RVT S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FADDX1_RVT S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FADDX1_RVT S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FADDX1_RVT S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FADDX1_RVT S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FADDX1_RVT S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FADDX1_RVT S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FADDX1_RVT S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FADDX1_RVT S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FADDX1_RVT S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FADDX1_RVT S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FADDX1_RVT S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FADDX1_RVT S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FADDX1_RVT S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FADDX1_RVT S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FADDX1_RVT S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FADDX1_RVT S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FADDX1_RVT S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FADDX1_RVT S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FADDX1_RVT S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FADDX1_RVT S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), 
        .CO(\CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FADDX1_RVT S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), 
        .CO(\CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FADDX1_RVT S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FADDX1_RVT S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FADDX1_RVT S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FADDX1_RVT S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), 
        .CO(\CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FADDX1_RVT S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), 
        .CO(\CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FADDX1_RVT S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), 
        .CO(\CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FADDX1_RVT S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), 
        .CO(\CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FADDX1_RVT S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FADDX1_RVT S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FADDX1_RVT S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FADDX1_RVT S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FADDX1_RVT S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), 
        .CO(\CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FADDX1_RVT S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), 
        .CO(\CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FADDX1_RVT S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), 
        .CO(\CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FADDX1_RVT S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FADDX1_RVT S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FADDX1_RVT S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), 
        .CO(\CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FADDX1_RVT S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), 
        .CO(\CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FADDX1_RVT S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), 
        .CO(\CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FADDX1_RVT S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), 
        .CO(\CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FADDX1_RVT S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), 
        .CO(\CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FADDX1_RVT S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), 
        .CO(\CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FADDX1_RVT S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), 
        .CO(\CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FADDX1_RVT S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), 
        .CO(\CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FADDX1_RVT S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), 
        .CO(\CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FADDX1_RVT S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FADDX1_RVT S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), 
        .CO(\CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FADDX1_RVT S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FADDX1_RVT S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), 
        .CO(\CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FADDX1_RVT S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FADDX1_RVT S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), 
        .CO(\CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FADDX1_RVT S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), 
        .CO(\CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FADDX1_RVT S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), 
        .CO(\CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FADDX1_RVT S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), 
        .CO(\CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FADDX1_RVT S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), 
        .CO(\CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FADDX1_RVT S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FADDX1_RVT S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), 
        .CO(\CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FADDX1_RVT S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), 
        .CO(\CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FADDX1_RVT S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FADDX1_RVT S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), 
        .CO(\CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FADDX1_RVT S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), 
        .CO(\CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FADDX1_RVT S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), 
        .CO(\CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FADDX1_RVT S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), 
        .CO(\CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FADDX1_RVT S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), 
        .CO(\CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FADDX1_RVT S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), 
        .CO(\CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FADDX1_RVT S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), 
        .CO(\CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FADDX1_RVT S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), 
        .CO(\CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FADDX1_RVT S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FADDX1_RVT S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), 
        .CO(\CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FADDX1_RVT S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), 
        .CO(\CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FADDX1_RVT S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), 
        .CO(\CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FADDX1_RVT S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), 
        .CO(\CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FADDX1_RVT S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FADDX1_RVT S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), 
        .CO(\CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FADDX1_RVT S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FADDX1_RVT S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FADDX1_RVT S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FADDX1_RVT S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), 
        .CO(\CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FADDX1_RVT S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), 
        .CO(\CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FADDX1_RVT S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), 
        .CO(\CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FADDX1_RVT S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), 
        .CO(\CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FADDX1_RVT S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), 
        .CO(\CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FADDX1_RVT S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FADDX1_RVT S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FADDX1_RVT S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FADDX1_RVT S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), 
        .CO(\CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FADDX1_RVT S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), 
        .CO(\CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FADDX1_RVT S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), 
        .CO(\CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FADDX1_RVT S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), 
        .CO(\CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FADDX1_RVT S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), 
        .CO(\CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FADDX1_RVT S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FADDX1_RVT S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), 
        .CO(\CARRYB[2][0] ), .S(\A1[0] ) );
  FADDX1_RVT S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), 
        .CO(\CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FADDX1_RVT S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), 
        .CO(\CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FADDX1_RVT S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), 
        .CO(\CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FADDX1_RVT S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), 
        .CO(\CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FADDX1_RVT S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), 
        .CO(\CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FADDX1_RVT S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), 
        .CO(\CARRYB[6][0] ), .S(\A1[4] ) );
  FADDX1_RVT S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), 
        .CO(\CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FADDX1_RVT S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), 
        .CO(\CARRYB[4][0] ), .S(\A1[2] ) );
  FADDX1_RVT S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), 
        .CO(\CARRYB[5][0] ), .S(\A1[3] ) );
  FADDX1_RVT S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), 
        .CO(\CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FADDX1_RVT S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), 
        .CO(\CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FADDX1_RVT S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), 
        .CO(\CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FADDX1_RVT S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), 
        .CO(\CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FADDX1_RVT S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FADDX1_RVT S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FADDX1_RVT S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FADDX1_RVT S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), 
        .CO(\CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FADDX1_RVT S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), 
        .CO(\CARRYB[8][0] ), .S(\A1[6] ) );
  FADDX1_RVT S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), 
        .CO(\CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FADDX1_RVT S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FADDX1_RVT S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), 
        .CO(\CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FADDX1_RVT S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FADDX1_RVT S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FADDX1_RVT S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), 
        .CO(\CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FADDX1_RVT S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), 
        .CO(\CARRYB[7][0] ), .S(\A1[5] ) );
  FADDX1_RVT S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), 
        .CO(\CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FADDX1_RVT S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), 
        .CO(\CARRYB[3][0] ), .S(\A1[1] ) );
  FADDX1_RVT S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), 
        .CO(\CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FADDX1_RVT S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), 
        .CO(\CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FADDX1_RVT S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), 
        .CO(\CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FADDX1_RVT S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), 
        .CO(\CARRYB[9][0] ), .S(\A1[7] ) );
  FADDX1_RVT S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), 
        .CO(\CARRYB[10][0] ), .S(\A1[8] ) );
  FADDX1_RVT S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FADDX1_RVT S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FADDX1_RVT S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FADDX1_RVT S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FADDX1_RVT S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FADDX1_RVT S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FADDX1_RVT S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FADDX1_RVT S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FADDX1_RVT S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FADDX1_RVT S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FADDX1_RVT S4_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FADDX1_RVT S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FADDX1_RVT S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FADDX1_RVT S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FADDX1_RVT S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), 
        .CO(\CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FADDX1_RVT S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), 
        .CO(\CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FADDX1_RVT S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), 
        .CO(\CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FADDX1_RVT S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), 
        .CO(\CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FADDX1_RVT S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), 
        .CO(\CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FADDX1_RVT S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), 
        .CO(\CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FADDX1_RVT S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FADDX1_RVT S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FADDX1_RVT S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FADDX1_RVT S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FADDX1_RVT S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), 
        .CO(\CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FADDX1_RVT S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), 
        .CO(\CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FADDX1_RVT S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), 
        .CO(\CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  IBUFFX2_RVT U2 ( .A(B[3]), .Y(n14) );
  INVX0_RVT U3 ( .A(B[23]), .Y(n74) );
  INVX0_RVT U4 ( .A(A[23]), .Y(n146) );
  INVX0_RVT U5 ( .A(A[21]), .Y(n140) );
  INVX0_RVT U6 ( .A(A[22]), .Y(n143) );
  INVX0_RVT U7 ( .A(B[22]), .Y(n71) );
  INVX0_RVT U8 ( .A(B[20]), .Y(n65) );
  INVX0_RVT U9 ( .A(B[21]), .Y(n68) );
  INVX0_RVT U10 ( .A(A[3]), .Y(n86) );
  INVX0_RVT U11 ( .A(A[5]), .Y(n92) );
  INVX0_RVT U12 ( .A(A[4]), .Y(n89) );
  INVX0_RVT U13 ( .A(A[6]), .Y(n95) );
  INVX0_RVT U14 ( .A(A[2]), .Y(n83) );
  INVX0_RVT U15 ( .A(A[1]), .Y(n80) );
  INVX0_RVT U16 ( .A(B[2]), .Y(n11) );
  INVX0_RVT U17 ( .A(A[8]), .Y(n101) );
  INVX0_RVT U18 ( .A(A[7]), .Y(n98) );
  INVX0_RVT U19 ( .A(A[9]), .Y(n104) );
  INVX0_RVT U20 ( .A(A[15]), .Y(n122) );
  INVX0_RVT U21 ( .A(A[13]), .Y(n116) );
  INVX0_RVT U22 ( .A(A[11]), .Y(n110) );
  INVX0_RVT U23 ( .A(A[17]), .Y(n128) );
  INVX0_RVT U24 ( .A(A[19]), .Y(n134) );
  INVX0_RVT U25 ( .A(A[16]), .Y(n125) );
  INVX0_RVT U26 ( .A(A[14]), .Y(n119) );
  INVX0_RVT U27 ( .A(A[12]), .Y(n113) );
  INVX0_RVT U28 ( .A(A[10]), .Y(n107) );
  INVX0_RVT U29 ( .A(A[18]), .Y(n131) );
  AND2X1_RVT U30 ( .A1(\ab[1][2] ), .A2(\ab[0][3] ), .Y(\CARRYB[1][2] ) );
  XOR2X1_RVT U31 ( .A1(\ab[0][4] ), .A2(\ab[1][3] ), .Y(\SUMB[1][3] ) );
  AND2X1_RVT U32 ( .A1(\CARRYB[23][2] ), .A2(\SUMB[23][3] ), .Y(\A2[25] ) );
  AND2X1_RVT U33 ( .A1(\CARRYB[23][5] ), .A2(\SUMB[23][6] ), .Y(\A2[28] ) );
  AND2X1_RVT U34 ( .A1(\CARRYB[23][6] ), .A2(\SUMB[23][7] ), .Y(\A2[29] ) );
  AND2X1_RVT U35 ( .A1(\CARRYB[23][7] ), .A2(\SUMB[23][8] ), .Y(\A2[30] ) );
  AND2X1_RVT U36 ( .A1(\CARRYB[23][8] ), .A2(\SUMB[23][9] ), .Y(\A2[31] ) );
  AND2X1_RVT U37 ( .A1(\CARRYB[23][9] ), .A2(\SUMB[23][10] ), .Y(\A2[32] ) );
  AND2X1_RVT U38 ( .A1(\CARRYB[23][1] ), .A2(\SUMB[23][2] ), .Y(\A2[24] ) );
  AND2X1_RVT U39 ( .A1(\CARRYB[23][3] ), .A2(\SUMB[23][4] ), .Y(\A2[26] ) );
  AND2X1_RVT U40 ( .A1(\CARRYB[23][0] ), .A2(\SUMB[23][1] ), .Y(\A2[23] ) );
  AND2X1_RVT U41 ( .A1(\CARRYB[23][4] ), .A2(\SUMB[23][5] ), .Y(\A2[27] ) );
  XOR2X1_RVT U42 ( .A1(\CARRYB[23][3] ), .A2(\SUMB[23][4] ), .Y(\A1[25] ) );
  XOR2X1_RVT U43 ( .A1(\CARRYB[23][6] ), .A2(\SUMB[23][7] ), .Y(\A1[28] ) );
  XOR2X1_RVT U44 ( .A1(\CARRYB[23][7] ), .A2(\SUMB[23][8] ), .Y(\A1[29] ) );
  XOR2X1_RVT U45 ( .A1(\CARRYB[23][8] ), .A2(\SUMB[23][9] ), .Y(\A1[30] ) );
  XOR2X1_RVT U46 ( .A1(\CARRYB[23][9] ), .A2(\SUMB[23][10] ), .Y(\A1[31] ) );
  XOR2X1_RVT U47 ( .A1(\CARRYB[23][10] ), .A2(\SUMB[23][11] ), .Y(\A1[32] ) );
  XOR2X1_RVT U48 ( .A1(\CARRYB[23][2] ), .A2(\SUMB[23][3] ), .Y(\A1[24] ) );
  XOR2X1_RVT U49 ( .A1(\CARRYB[23][4] ), .A2(\SUMB[23][5] ), .Y(\A1[26] ) );
  XOR2X1_RVT U50 ( .A1(\CARRYB[23][1] ), .A2(\SUMB[23][2] ), .Y(\A1[23] ) );
  XOR2X1_RVT U51 ( .A1(\CARRYB[23][5] ), .A2(\SUMB[23][6] ), .Y(\A1[27] ) );
  AND2X1_RVT U52 ( .A1(\CARRYB[23][21] ), .A2(\SUMB[23][22] ), .Y(\A2[44] ) );
  XOR2X1_RVT U53 ( .A1(\CARRYB[23][22] ), .A2(\ab[23][23] ), .Y(\A1[44] ) );
  AND2X1_RVT U54 ( .A1(\CARRYB[23][10] ), .A2(\SUMB[23][11] ), .Y(\A2[33] ) );
  AND2X1_RVT U55 ( .A1(\CARRYB[23][11] ), .A2(\SUMB[23][12] ), .Y(\A2[34] ) );
  AND2X1_RVT U56 ( .A1(\CARRYB[23][12] ), .A2(\SUMB[23][13] ), .Y(\A2[35] ) );
  AND2X1_RVT U57 ( .A1(\CARRYB[23][13] ), .A2(\SUMB[23][14] ), .Y(\A2[36] ) );
  AND2X1_RVT U58 ( .A1(\CARRYB[23][14] ), .A2(\SUMB[23][15] ), .Y(\A2[37] ) );
  AND2X1_RVT U59 ( .A1(\CARRYB[23][15] ), .A2(\SUMB[23][16] ), .Y(\A2[38] ) );
  AND2X1_RVT U60 ( .A1(\CARRYB[23][16] ), .A2(\SUMB[23][17] ), .Y(\A2[39] ) );
  AND2X1_RVT U61 ( .A1(\CARRYB[23][17] ), .A2(\SUMB[23][18] ), .Y(\A2[40] ) );
  AND2X1_RVT U62 ( .A1(\CARRYB[23][18] ), .A2(\SUMB[23][19] ), .Y(\A2[41] ) );
  AND2X1_RVT U63 ( .A1(\CARRYB[23][19] ), .A2(\SUMB[23][20] ), .Y(\A2[42] ) );
  AND2X1_RVT U64 ( .A1(\CARRYB[23][20] ), .A2(\SUMB[23][21] ), .Y(\A2[43] ) );
  XOR2X1_RVT U65 ( .A1(\CARRYB[23][11] ), .A2(\SUMB[23][12] ), .Y(\A1[33] ) );
  XOR2X1_RVT U66 ( .A1(\CARRYB[23][12] ), .A2(\SUMB[23][13] ), .Y(\A1[34] ) );
  XOR2X1_RVT U67 ( .A1(\CARRYB[23][13] ), .A2(\SUMB[23][14] ), .Y(\A1[35] ) );
  XOR2X1_RVT U68 ( .A1(\CARRYB[23][14] ), .A2(\SUMB[23][15] ), .Y(\A1[36] ) );
  XOR2X1_RVT U69 ( .A1(\CARRYB[23][15] ), .A2(\SUMB[23][16] ), .Y(\A1[37] ) );
  XOR2X1_RVT U70 ( .A1(\CARRYB[23][16] ), .A2(\SUMB[23][17] ), .Y(\A1[38] ) );
  XOR2X1_RVT U71 ( .A1(\CARRYB[23][17] ), .A2(\SUMB[23][18] ), .Y(\A1[39] ) );
  XOR2X1_RVT U72 ( .A1(\CARRYB[23][18] ), .A2(\SUMB[23][19] ), .Y(\A1[40] ) );
  XOR2X1_RVT U73 ( .A1(\CARRYB[23][19] ), .A2(\SUMB[23][20] ), .Y(\A1[41] ) );
  XOR2X1_RVT U74 ( .A1(\CARRYB[23][20] ), .A2(\SUMB[23][21] ), .Y(\A1[42] ) );
  XOR2X1_RVT U75 ( .A1(\CARRYB[23][21] ), .A2(\SUMB[23][22] ), .Y(\A1[43] ) );
  XOR2X1_RVT U76 ( .A1(\ab[0][1] ), .A2(\ab[1][0] ), .Y(PRODUCT[1]) );
  INVX1_RVT U77 ( .A(n104), .Y(n102) );
  INVX1_RVT U78 ( .A(n104), .Y(n103) );
  INVX1_RVT U79 ( .A(n86), .Y(n84) );
  INVX1_RVT U80 ( .A(n86), .Y(n85) );
  INVX1_RVT U81 ( .A(n98), .Y(n96) );
  INVX1_RVT U82 ( .A(n98), .Y(n97) );
  INVX1_RVT U83 ( .A(n110), .Y(n109) );
  INVX1_RVT U84 ( .A(n101), .Y(n99) );
  INVX1_RVT U85 ( .A(n113), .Y(n112) );
  INVX1_RVT U86 ( .A(n101), .Y(n100) );
  INVX1_RVT U87 ( .A(n107), .Y(n106) );
  INVX1_RVT U88 ( .A(n107), .Y(n105) );
  INVX1_RVT U89 ( .A(n92), .Y(n90) );
  INVX1_RVT U90 ( .A(n92), .Y(n91) );
  INVX1_RVT U91 ( .A(n89), .Y(n87) );
  INVX1_RVT U92 ( .A(n95), .Y(n93) );
  INVX1_RVT U93 ( .A(n89), .Y(n88) );
  INVX1_RVT U94 ( .A(n95), .Y(n94) );
  INVX1_RVT U95 ( .A(n80), .Y(n78) );
  INVX1_RVT U96 ( .A(n80), .Y(n79) );
  INVX1_RVT U97 ( .A(n11), .Y(n10) );
  INVX1_RVT U98 ( .A(n77), .Y(n76) );
  INVX1_RVT U99 ( .A(n77), .Y(n75) );
  INVX1_RVT U100 ( .A(n83), .Y(n81) );
  INVX1_RVT U101 ( .A(n83), .Y(n82) );
  INVX1_RVT U102 ( .A(n11), .Y(n9) );
  XOR2X1_RVT U103 ( .A1(\ab[0][3] ), .A2(\ab[1][2] ), .Y(\SUMB[1][2] ) );
  AND2X1_RVT U104 ( .A1(\ab[1][1] ), .A2(\ab[0][2] ), .Y(\CARRYB[1][1] ) );
  XOR2X1_RVT U105 ( .A1(\ab[0][2] ), .A2(\ab[1][1] ), .Y(\SUMB[1][1] ) );
  AND2X1_RVT U106 ( .A1(\ab[1][0] ), .A2(\ab[0][1] ), .Y(\CARRYB[1][0] ) );
  XOR2X1_RVT U107 ( .A1(\ab[0][5] ), .A2(\ab[1][4] ), .Y(\SUMB[1][4] ) );
  AND2X1_RVT U108 ( .A1(\ab[1][3] ), .A2(\ab[0][4] ), .Y(\CARRYB[1][3] ) );
  AND2X1_RVT U109 ( .A1(\ab[1][4] ), .A2(\ab[0][5] ), .Y(\CARRYB[1][4] ) );
  XOR2X1_RVT U110 ( .A1(\ab[0][6] ), .A2(\ab[1][5] ), .Y(\SUMB[1][5] ) );
  XOR2X1_RVT U111 ( .A1(\ab[0][7] ), .A2(\ab[1][6] ), .Y(\SUMB[1][6] ) );
  AND2X1_RVT U112 ( .A1(\ab[1][5] ), .A2(\ab[0][6] ), .Y(\CARRYB[1][5] ) );
  XOR2X1_RVT U113 ( .A1(\ab[0][15] ), .A2(\ab[1][14] ), .Y(\SUMB[1][14] ) );
  AND2X1_RVT U114 ( .A1(\ab[1][13] ), .A2(\ab[0][14] ), .Y(\CARRYB[1][13] ) );
  AND2X1_RVT U115 ( .A1(\ab[1][12] ), .A2(\ab[0][13] ), .Y(\CARRYB[1][12] ) );
  XOR2X1_RVT U116 ( .A1(\ab[0][14] ), .A2(\ab[1][13] ), .Y(\SUMB[1][13] ) );
  XOR2X1_RVT U117 ( .A1(\ab[0][13] ), .A2(\ab[1][12] ), .Y(\SUMB[1][12] ) );
  AND2X1_RVT U118 ( .A1(\ab[1][11] ), .A2(\ab[0][12] ), .Y(\CARRYB[1][11] ) );
  AND2X1_RVT U119 ( .A1(\ab[1][10] ), .A2(\ab[0][11] ), .Y(\CARRYB[1][10] ) );
  XOR2X1_RVT U120 ( .A1(\ab[0][12] ), .A2(\ab[1][11] ), .Y(\SUMB[1][11] ) );
  XOR2X1_RVT U121 ( .A1(\ab[0][11] ), .A2(\ab[1][10] ), .Y(\SUMB[1][10] ) );
  AND2X1_RVT U122 ( .A1(\ab[1][9] ), .A2(\ab[0][10] ), .Y(\CARRYB[1][9] ) );
  AND2X1_RVT U123 ( .A1(\ab[1][8] ), .A2(\ab[0][9] ), .Y(\CARRYB[1][8] ) );
  XOR2X1_RVT U124 ( .A1(\ab[0][10] ), .A2(\ab[1][9] ), .Y(\SUMB[1][9] ) );
  XOR2X1_RVT U125 ( .A1(\ab[0][9] ), .A2(\ab[1][8] ), .Y(\SUMB[1][8] ) );
  AND2X1_RVT U126 ( .A1(\ab[1][7] ), .A2(\ab[0][8] ), .Y(\CARRYB[1][7] ) );
  AND2X1_RVT U127 ( .A1(\ab[1][6] ), .A2(\ab[0][7] ), .Y(\CARRYB[1][6] ) );
  XOR2X1_RVT U128 ( .A1(\ab[0][8] ), .A2(\ab[1][7] ), .Y(\SUMB[1][7] ) );
  AND2X1_RVT U129 ( .A1(\ab[1][14] ), .A2(\ab[0][15] ), .Y(\CARRYB[1][14] ) );
  XOR2X1_RVT U130 ( .A1(\ab[0][16] ), .A2(\ab[1][15] ), .Y(\SUMB[1][15] ) );
  INVX1_RVT U131 ( .A(n125), .Y(n123) );
  INVX1_RVT U132 ( .A(n122), .Y(n120) );
  INVX1_RVT U133 ( .A(n116), .Y(n115) );
  INVX1_RVT U134 ( .A(n116), .Y(n114) );
  INVX1_RVT U135 ( .A(n110), .Y(n108) );
  INVX1_RVT U136 ( .A(n119), .Y(n117) );
  INVX1_RVT U137 ( .A(n119), .Y(n118) );
  INVX1_RVT U138 ( .A(n113), .Y(n111) );
  AND2X1_RVT U139 ( .A1(\ab[1][16] ), .A2(\ab[0][17] ), .Y(\CARRYB[1][16] ) );
  XOR2X1_RVT U140 ( .A1(\ab[0][18] ), .A2(\ab[1][17] ), .Y(\SUMB[1][17] ) );
  AND2X1_RVT U141 ( .A1(\ab[1][15] ), .A2(\ab[0][16] ), .Y(\CARRYB[1][15] ) );
  XOR2X1_RVT U142 ( .A1(\ab[0][17] ), .A2(\ab[1][16] ), .Y(\SUMB[1][16] ) );
  AND2X1_RVT U143 ( .A1(\ab[1][17] ), .A2(\ab[0][18] ), .Y(\CARRYB[1][17] ) );
  XOR2X1_RVT U144 ( .A1(\ab[0][19] ), .A2(\ab[1][18] ), .Y(\SUMB[1][18] ) );
  INVX1_RVT U145 ( .A(n128), .Y(n127) );
  INVX1_RVT U146 ( .A(n128), .Y(n126) );
  INVX1_RVT U147 ( .A(n134), .Y(n132) );
  INVX1_RVT U148 ( .A(n125), .Y(n124) );
  INVX1_RVT U149 ( .A(n131), .Y(n129) );
  INVX1_RVT U150 ( .A(n122), .Y(n121) );
  AND2X1_RVT U151 ( .A1(\CARRYB[23][22] ), .A2(\ab[23][23] ), .Y(\A2[45] ) );
  INVX1_RVT U152 ( .A(n74), .Y(n73) );
  INVX1_RVT U153 ( .A(n74), .Y(n72) );
  AND2X1_RVT U154 ( .A1(\ab[1][22] ), .A2(\ab[0][23] ), .Y(\CARRYB[1][22] ) );
  AND2X1_RVT U155 ( .A1(\ab[1][21] ), .A2(\ab[0][22] ), .Y(\CARRYB[1][21] ) );
  XOR2X1_RVT U156 ( .A1(\ab[0][23] ), .A2(\ab[1][22] ), .Y(\SUMB[1][22] ) );
  AND2X1_RVT U157 ( .A1(\ab[1][20] ), .A2(\ab[0][21] ), .Y(\CARRYB[1][20] ) );
  XOR2X1_RVT U158 ( .A1(\ab[0][22] ), .A2(\ab[1][21] ), .Y(\SUMB[1][21] ) );
  AND2X1_RVT U159 ( .A1(\ab[1][19] ), .A2(\ab[0][20] ), .Y(\CARRYB[1][19] ) );
  XOR2X1_RVT U160 ( .A1(\ab[0][21] ), .A2(\ab[1][20] ), .Y(\SUMB[1][20] ) );
  AND2X1_RVT U161 ( .A1(\ab[1][18] ), .A2(\ab[0][19] ), .Y(\CARRYB[1][18] ) );
  XOR2X1_RVT U162 ( .A1(\ab[0][20] ), .A2(\ab[1][19] ), .Y(\SUMB[1][19] ) );
  INVX1_RVT U163 ( .A(n140), .Y(n139) );
  INVX1_RVT U164 ( .A(n140), .Y(n138) );
  INVX1_RVT U165 ( .A(n134), .Y(n133) );
  INVX1_RVT U166 ( .A(n131), .Y(n130) );
  INVX1_RVT U167 ( .A(n137), .Y(n136) );
  INVX1_RVT U168 ( .A(n137), .Y(n135) );
  INVX1_RVT U169 ( .A(n143), .Y(n142) );
  INVX1_RVT U170 ( .A(n143), .Y(n141) );
  INVX1_RVT U171 ( .A(n146), .Y(n145) );
  INVX1_RVT U172 ( .A(n146), .Y(n144) );
  XOR2X1_RVT U173 ( .A1(\CARRYB[23][0] ), .A2(\SUMB[23][1] ), .Y(\A1[22] ) );
  INVX1_RVT U174 ( .A(n5), .Y(n3) );
  INVX1_RVT U175 ( .A(A[0]), .Y(n77) );
  INVX1_RVT U176 ( .A(n8), .Y(n6) );
  INVX1_RVT U177 ( .A(n14), .Y(n12) );
  INVX1_RVT U178 ( .A(n17), .Y(n15) );
  INVX1_RVT U179 ( .A(n50), .Y(n48) );
  INVX1_RVT U180 ( .A(n47), .Y(n45) );
  INVX1_RVT U181 ( .A(n44), .Y(n42) );
  INVX1_RVT U182 ( .A(n41), .Y(n39) );
  INVX1_RVT U183 ( .A(n38), .Y(n36) );
  INVX1_RVT U184 ( .A(n35), .Y(n33) );
  INVX1_RVT U185 ( .A(n32), .Y(n30) );
  INVX1_RVT U186 ( .A(n29), .Y(n27) );
  INVX1_RVT U187 ( .A(n26), .Y(n24) );
  INVX1_RVT U188 ( .A(n23), .Y(n21) );
  INVX1_RVT U189 ( .A(n20), .Y(n18) );
  INVX1_RVT U190 ( .A(n8), .Y(n7) );
  INVX1_RVT U191 ( .A(n14), .Y(n13) );
  INVX1_RVT U192 ( .A(n17), .Y(n16) );
  INVX1_RVT U193 ( .A(n50), .Y(n49) );
  INVX1_RVT U194 ( .A(n53), .Y(n52) );
  INVX1_RVT U195 ( .A(n47), .Y(n46) );
  INVX1_RVT U196 ( .A(n44), .Y(n43) );
  INVX1_RVT U197 ( .A(n38), .Y(n37) );
  INVX1_RVT U198 ( .A(n41), .Y(n40) );
  INVX1_RVT U199 ( .A(n32), .Y(n31) );
  INVX1_RVT U200 ( .A(n35), .Y(n34) );
  INVX1_RVT U201 ( .A(n20), .Y(n19) );
  INVX1_RVT U202 ( .A(n29), .Y(n28) );
  INVX1_RVT U203 ( .A(n26), .Y(n25) );
  INVX1_RVT U204 ( .A(n23), .Y(n22) );
  INVX1_RVT U205 ( .A(n5), .Y(n4) );
  INVX1_RVT U206 ( .A(n59), .Y(n57) );
  INVX1_RVT U207 ( .A(n56), .Y(n54) );
  INVX1_RVT U208 ( .A(n53), .Y(n51) );
  INVX1_RVT U209 ( .A(n59), .Y(n58) );
  INVX1_RVT U210 ( .A(n62), .Y(n61) );
  INVX1_RVT U211 ( .A(n56), .Y(n55) );
  INVX1_RVT U212 ( .A(n65), .Y(n63) );
  INVX1_RVT U213 ( .A(n62), .Y(n60) );
  INVX1_RVT U214 ( .A(n68), .Y(n66) );
  INVX1_RVT U215 ( .A(n71), .Y(n69) );
  INVX1_RVT U216 ( .A(n71), .Y(n70) );
  INVX1_RVT U217 ( .A(n68), .Y(n67) );
  INVX1_RVT U218 ( .A(n65), .Y(n64) );
  INVX1_RVT U219 ( .A(A[20]), .Y(n137) );
  INVX1_RVT U220 ( .A(B[9]), .Y(n32) );
  INVX1_RVT U221 ( .A(B[7]), .Y(n26) );
  INVX1_RVT U222 ( .A(B[15]), .Y(n50) );
  INVX1_RVT U223 ( .A(B[5]), .Y(n20) );
  INVX1_RVT U224 ( .A(B[4]), .Y(n17) );
  INVX1_RVT U225 ( .A(B[13]), .Y(n44) );
  INVX1_RVT U226 ( .A(B[11]), .Y(n38) );
  INVX1_RVT U227 ( .A(B[8]), .Y(n29) );
  INVX1_RVT U228 ( .A(B[6]), .Y(n23) );
  INVX1_RVT U229 ( .A(B[14]), .Y(n47) );
  INVX1_RVT U230 ( .A(B[12]), .Y(n41) );
  INVX1_RVT U231 ( .A(B[10]), .Y(n35) );
  INVX1_RVT U232 ( .A(B[16]), .Y(n53) );
  INVX1_RVT U233 ( .A(B[1]), .Y(n8) );
  INVX1_RVT U234 ( .A(B[0]), .Y(n5) );
  INVX1_RVT U235 ( .A(B[19]), .Y(n62) );
  INVX1_RVT U236 ( .A(B[17]), .Y(n56) );
  INVX1_RVT U237 ( .A(B[18]), .Y(n59) );
  AND2X1_RVT U239 ( .A1(n30), .A2(n103), .Y(\ab[9][9] ) );
  AND2X1_RVT U240 ( .A1(n27), .A2(n103), .Y(\ab[9][8] ) );
  AND2X1_RVT U241 ( .A1(n24), .A2(n103), .Y(\ab[9][7] ) );
  AND2X1_RVT U242 ( .A1(n21), .A2(n103), .Y(\ab[9][6] ) );
  AND2X1_RVT U243 ( .A1(n18), .A2(n103), .Y(\ab[9][5] ) );
  AND2X1_RVT U244 ( .A1(n15), .A2(n103), .Y(\ab[9][4] ) );
  AND2X1_RVT U245 ( .A1(n12), .A2(n103), .Y(\ab[9][3] ) );
  AND2X1_RVT U246 ( .A1(n9), .A2(n103), .Y(\ab[9][2] ) );
  AND2X1_RVT U247 ( .A1(n72), .A2(n103), .Y(\ab[9][23] ) );
  AND2X1_RVT U248 ( .A1(n69), .A2(n103), .Y(\ab[9][22] ) );
  AND2X1_RVT U249 ( .A1(n66), .A2(n103), .Y(\ab[9][21] ) );
  AND2X1_RVT U250 ( .A1(n63), .A2(n103), .Y(\ab[9][20] ) );
  AND2X1_RVT U251 ( .A1(n6), .A2(n102), .Y(\ab[9][1] ) );
  AND2X1_RVT U252 ( .A1(n60), .A2(n102), .Y(\ab[9][19] ) );
  AND2X1_RVT U253 ( .A1(n57), .A2(n102), .Y(\ab[9][18] ) );
  AND2X1_RVT U254 ( .A1(n54), .A2(n102), .Y(\ab[9][17] ) );
  AND2X1_RVT U255 ( .A1(n51), .A2(n102), .Y(\ab[9][16] ) );
  AND2X1_RVT U256 ( .A1(n48), .A2(n102), .Y(\ab[9][15] ) );
  AND2X1_RVT U257 ( .A1(n45), .A2(n102), .Y(\ab[9][14] ) );
  AND2X1_RVT U258 ( .A1(n42), .A2(n102), .Y(\ab[9][13] ) );
  AND2X1_RVT U259 ( .A1(n39), .A2(n102), .Y(\ab[9][12] ) );
  AND2X1_RVT U260 ( .A1(n36), .A2(n102), .Y(\ab[9][11] ) );
  AND2X1_RVT U261 ( .A1(n33), .A2(n102), .Y(\ab[9][10] ) );
  AND2X1_RVT U262 ( .A1(n3), .A2(n102), .Y(\ab[9][0] ) );
  AND2X1_RVT U263 ( .A1(n100), .A2(n30), .Y(\ab[8][9] ) );
  AND2X1_RVT U264 ( .A1(n100), .A2(n27), .Y(\ab[8][8] ) );
  AND2X1_RVT U265 ( .A1(n100), .A2(n24), .Y(\ab[8][7] ) );
  AND2X1_RVT U266 ( .A1(n100), .A2(n21), .Y(\ab[8][6] ) );
  AND2X1_RVT U267 ( .A1(n100), .A2(n18), .Y(\ab[8][5] ) );
  AND2X1_RVT U268 ( .A1(n100), .A2(n15), .Y(\ab[8][4] ) );
  AND2X1_RVT U269 ( .A1(n100), .A2(n12), .Y(\ab[8][3] ) );
  AND2X1_RVT U270 ( .A1(n100), .A2(n9), .Y(\ab[8][2] ) );
  AND2X1_RVT U271 ( .A1(n100), .A2(n72), .Y(\ab[8][23] ) );
  AND2X1_RVT U272 ( .A1(n100), .A2(n69), .Y(\ab[8][22] ) );
  AND2X1_RVT U273 ( .A1(n100), .A2(n66), .Y(\ab[8][21] ) );
  AND2X1_RVT U274 ( .A1(n100), .A2(n63), .Y(\ab[8][20] ) );
  AND2X1_RVT U275 ( .A1(n99), .A2(n6), .Y(\ab[8][1] ) );
  AND2X1_RVT U276 ( .A1(n99), .A2(n60), .Y(\ab[8][19] ) );
  AND2X1_RVT U277 ( .A1(n99), .A2(n57), .Y(\ab[8][18] ) );
  AND2X1_RVT U278 ( .A1(n99), .A2(n54), .Y(\ab[8][17] ) );
  AND2X1_RVT U279 ( .A1(n99), .A2(n51), .Y(\ab[8][16] ) );
  AND2X1_RVT U280 ( .A1(n99), .A2(n48), .Y(\ab[8][15] ) );
  AND2X1_RVT U281 ( .A1(n99), .A2(n45), .Y(\ab[8][14] ) );
  AND2X1_RVT U282 ( .A1(n99), .A2(n42), .Y(\ab[8][13] ) );
  AND2X1_RVT U283 ( .A1(n99), .A2(n39), .Y(\ab[8][12] ) );
  AND2X1_RVT U284 ( .A1(n99), .A2(n36), .Y(\ab[8][11] ) );
  AND2X1_RVT U285 ( .A1(n99), .A2(n33), .Y(\ab[8][10] ) );
  AND2X1_RVT U286 ( .A1(n99), .A2(n3), .Y(\ab[8][0] ) );
  AND2X1_RVT U287 ( .A1(n97), .A2(n30), .Y(\ab[7][9] ) );
  AND2X1_RVT U288 ( .A1(n97), .A2(n27), .Y(\ab[7][8] ) );
  AND2X1_RVT U289 ( .A1(n97), .A2(n24), .Y(\ab[7][7] ) );
  AND2X1_RVT U290 ( .A1(n97), .A2(n21), .Y(\ab[7][6] ) );
  AND2X1_RVT U291 ( .A1(n97), .A2(n18), .Y(\ab[7][5] ) );
  AND2X1_RVT U292 ( .A1(n97), .A2(n15), .Y(\ab[7][4] ) );
  AND2X1_RVT U293 ( .A1(n97), .A2(n12), .Y(\ab[7][3] ) );
  AND2X1_RVT U294 ( .A1(n97), .A2(n9), .Y(\ab[7][2] ) );
  AND2X1_RVT U295 ( .A1(n97), .A2(n72), .Y(\ab[7][23] ) );
  AND2X1_RVT U296 ( .A1(n97), .A2(n69), .Y(\ab[7][22] ) );
  AND2X1_RVT U297 ( .A1(n97), .A2(n66), .Y(\ab[7][21] ) );
  AND2X1_RVT U298 ( .A1(n97), .A2(n63), .Y(\ab[7][20] ) );
  AND2X1_RVT U299 ( .A1(n96), .A2(n6), .Y(\ab[7][1] ) );
  AND2X1_RVT U300 ( .A1(n96), .A2(n60), .Y(\ab[7][19] ) );
  AND2X1_RVT U301 ( .A1(n96), .A2(n57), .Y(\ab[7][18] ) );
  AND2X1_RVT U302 ( .A1(n96), .A2(n54), .Y(\ab[7][17] ) );
  AND2X1_RVT U303 ( .A1(n96), .A2(n51), .Y(\ab[7][16] ) );
  AND2X1_RVT U304 ( .A1(n96), .A2(n48), .Y(\ab[7][15] ) );
  AND2X1_RVT U305 ( .A1(n96), .A2(n45), .Y(\ab[7][14] ) );
  AND2X1_RVT U306 ( .A1(n96), .A2(n42), .Y(\ab[7][13] ) );
  AND2X1_RVT U307 ( .A1(n96), .A2(n39), .Y(\ab[7][12] ) );
  AND2X1_RVT U308 ( .A1(n96), .A2(n36), .Y(\ab[7][11] ) );
  AND2X1_RVT U309 ( .A1(n96), .A2(n33), .Y(\ab[7][10] ) );
  AND2X1_RVT U310 ( .A1(n96), .A2(n3), .Y(\ab[7][0] ) );
  AND2X1_RVT U311 ( .A1(n94), .A2(n30), .Y(\ab[6][9] ) );
  AND2X1_RVT U312 ( .A1(n94), .A2(n27), .Y(\ab[6][8] ) );
  AND2X1_RVT U313 ( .A1(n94), .A2(n24), .Y(\ab[6][7] ) );
  AND2X1_RVT U314 ( .A1(n94), .A2(n21), .Y(\ab[6][6] ) );
  AND2X1_RVT U315 ( .A1(n94), .A2(n18), .Y(\ab[6][5] ) );
  AND2X1_RVT U316 ( .A1(n94), .A2(n15), .Y(\ab[6][4] ) );
  AND2X1_RVT U317 ( .A1(n94), .A2(n12), .Y(\ab[6][3] ) );
  AND2X1_RVT U318 ( .A1(n94), .A2(n9), .Y(\ab[6][2] ) );
  AND2X1_RVT U319 ( .A1(n94), .A2(n72), .Y(\ab[6][23] ) );
  AND2X1_RVT U320 ( .A1(n94), .A2(n69), .Y(\ab[6][22] ) );
  AND2X1_RVT U321 ( .A1(n94), .A2(n66), .Y(\ab[6][21] ) );
  AND2X1_RVT U322 ( .A1(n94), .A2(n63), .Y(\ab[6][20] ) );
  AND2X1_RVT U323 ( .A1(n93), .A2(n6), .Y(\ab[6][1] ) );
  AND2X1_RVT U324 ( .A1(n93), .A2(n60), .Y(\ab[6][19] ) );
  AND2X1_RVT U325 ( .A1(n93), .A2(n57), .Y(\ab[6][18] ) );
  AND2X1_RVT U326 ( .A1(n93), .A2(n54), .Y(\ab[6][17] ) );
  AND2X1_RVT U327 ( .A1(n93), .A2(n51), .Y(\ab[6][16] ) );
  AND2X1_RVT U328 ( .A1(n93), .A2(n48), .Y(\ab[6][15] ) );
  AND2X1_RVT U329 ( .A1(n93), .A2(n45), .Y(\ab[6][14] ) );
  AND2X1_RVT U330 ( .A1(n93), .A2(n42), .Y(\ab[6][13] ) );
  AND2X1_RVT U331 ( .A1(n93), .A2(n39), .Y(\ab[6][12] ) );
  AND2X1_RVT U332 ( .A1(n93), .A2(n36), .Y(\ab[6][11] ) );
  AND2X1_RVT U333 ( .A1(n93), .A2(n33), .Y(\ab[6][10] ) );
  AND2X1_RVT U334 ( .A1(n93), .A2(n3), .Y(\ab[6][0] ) );
  AND2X1_RVT U335 ( .A1(n91), .A2(n30), .Y(\ab[5][9] ) );
  AND2X1_RVT U336 ( .A1(n91), .A2(n27), .Y(\ab[5][8] ) );
  AND2X1_RVT U337 ( .A1(n91), .A2(n24), .Y(\ab[5][7] ) );
  AND2X1_RVT U338 ( .A1(n91), .A2(n21), .Y(\ab[5][6] ) );
  AND2X1_RVT U339 ( .A1(n91), .A2(n18), .Y(\ab[5][5] ) );
  AND2X1_RVT U340 ( .A1(n91), .A2(n15), .Y(\ab[5][4] ) );
  AND2X1_RVT U341 ( .A1(n91), .A2(n12), .Y(\ab[5][3] ) );
  AND2X1_RVT U342 ( .A1(n91), .A2(n9), .Y(\ab[5][2] ) );
  AND2X1_RVT U343 ( .A1(n91), .A2(n72), .Y(\ab[5][23] ) );
  AND2X1_RVT U344 ( .A1(n91), .A2(n69), .Y(\ab[5][22] ) );
  AND2X1_RVT U345 ( .A1(n91), .A2(n66), .Y(\ab[5][21] ) );
  AND2X1_RVT U346 ( .A1(n91), .A2(n63), .Y(\ab[5][20] ) );
  AND2X1_RVT U347 ( .A1(n90), .A2(n6), .Y(\ab[5][1] ) );
  AND2X1_RVT U348 ( .A1(n90), .A2(n60), .Y(\ab[5][19] ) );
  AND2X1_RVT U349 ( .A1(n90), .A2(n57), .Y(\ab[5][18] ) );
  AND2X1_RVT U350 ( .A1(n90), .A2(n54), .Y(\ab[5][17] ) );
  AND2X1_RVT U351 ( .A1(n90), .A2(n51), .Y(\ab[5][16] ) );
  AND2X1_RVT U352 ( .A1(n90), .A2(n48), .Y(\ab[5][15] ) );
  AND2X1_RVT U353 ( .A1(n90), .A2(n45), .Y(\ab[5][14] ) );
  AND2X1_RVT U354 ( .A1(n90), .A2(n42), .Y(\ab[5][13] ) );
  AND2X1_RVT U355 ( .A1(n90), .A2(n39), .Y(\ab[5][12] ) );
  AND2X1_RVT U356 ( .A1(n90), .A2(n36), .Y(\ab[5][11] ) );
  AND2X1_RVT U357 ( .A1(n90), .A2(n33), .Y(\ab[5][10] ) );
  AND2X1_RVT U358 ( .A1(n90), .A2(n3), .Y(\ab[5][0] ) );
  AND2X1_RVT U359 ( .A1(n88), .A2(n30), .Y(\ab[4][9] ) );
  AND2X1_RVT U360 ( .A1(n88), .A2(n27), .Y(\ab[4][8] ) );
  AND2X1_RVT U361 ( .A1(n88), .A2(n24), .Y(\ab[4][7] ) );
  AND2X1_RVT U362 ( .A1(n88), .A2(n21), .Y(\ab[4][6] ) );
  AND2X1_RVT U363 ( .A1(n88), .A2(n18), .Y(\ab[4][5] ) );
  AND2X1_RVT U364 ( .A1(n88), .A2(n15), .Y(\ab[4][4] ) );
  AND2X1_RVT U365 ( .A1(n88), .A2(n12), .Y(\ab[4][3] ) );
  AND2X1_RVT U366 ( .A1(n88), .A2(n9), .Y(\ab[4][2] ) );
  AND2X1_RVT U367 ( .A1(n88), .A2(n72), .Y(\ab[4][23] ) );
  AND2X1_RVT U368 ( .A1(n88), .A2(n69), .Y(\ab[4][22] ) );
  AND2X1_RVT U369 ( .A1(n88), .A2(n66), .Y(\ab[4][21] ) );
  AND2X1_RVT U370 ( .A1(n88), .A2(n63), .Y(\ab[4][20] ) );
  AND2X1_RVT U371 ( .A1(n87), .A2(n6), .Y(\ab[4][1] ) );
  AND2X1_RVT U372 ( .A1(n87), .A2(n60), .Y(\ab[4][19] ) );
  AND2X1_RVT U373 ( .A1(n87), .A2(n57), .Y(\ab[4][18] ) );
  AND2X1_RVT U374 ( .A1(n87), .A2(n54), .Y(\ab[4][17] ) );
  AND2X1_RVT U375 ( .A1(n87), .A2(n51), .Y(\ab[4][16] ) );
  AND2X1_RVT U376 ( .A1(n87), .A2(n48), .Y(\ab[4][15] ) );
  AND2X1_RVT U377 ( .A1(n87), .A2(n45), .Y(\ab[4][14] ) );
  AND2X1_RVT U378 ( .A1(n87), .A2(n42), .Y(\ab[4][13] ) );
  AND2X1_RVT U379 ( .A1(n87), .A2(n39), .Y(\ab[4][12] ) );
  AND2X1_RVT U380 ( .A1(n87), .A2(n36), .Y(\ab[4][11] ) );
  AND2X1_RVT U381 ( .A1(n87), .A2(n33), .Y(\ab[4][10] ) );
  AND2X1_RVT U382 ( .A1(n87), .A2(n3), .Y(\ab[4][0] ) );
  AND2X1_RVT U383 ( .A1(n85), .A2(n30), .Y(\ab[3][9] ) );
  AND2X1_RVT U384 ( .A1(n85), .A2(n27), .Y(\ab[3][8] ) );
  AND2X1_RVT U385 ( .A1(n85), .A2(n24), .Y(\ab[3][7] ) );
  AND2X1_RVT U386 ( .A1(n85), .A2(n21), .Y(\ab[3][6] ) );
  AND2X1_RVT U387 ( .A1(n85), .A2(n18), .Y(\ab[3][5] ) );
  AND2X1_RVT U388 ( .A1(n85), .A2(n15), .Y(\ab[3][4] ) );
  AND2X1_RVT U389 ( .A1(n85), .A2(n12), .Y(\ab[3][3] ) );
  AND2X1_RVT U390 ( .A1(n85), .A2(n9), .Y(\ab[3][2] ) );
  AND2X1_RVT U391 ( .A1(n85), .A2(n72), .Y(\ab[3][23] ) );
  AND2X1_RVT U392 ( .A1(n85), .A2(n69), .Y(\ab[3][22] ) );
  AND2X1_RVT U393 ( .A1(n85), .A2(n66), .Y(\ab[3][21] ) );
  AND2X1_RVT U394 ( .A1(n85), .A2(n63), .Y(\ab[3][20] ) );
  AND2X1_RVT U395 ( .A1(n84), .A2(n6), .Y(\ab[3][1] ) );
  AND2X1_RVT U396 ( .A1(n84), .A2(n60), .Y(\ab[3][19] ) );
  AND2X1_RVT U397 ( .A1(n84), .A2(n57), .Y(\ab[3][18] ) );
  AND2X1_RVT U398 ( .A1(n84), .A2(n54), .Y(\ab[3][17] ) );
  AND2X1_RVT U399 ( .A1(n84), .A2(n51), .Y(\ab[3][16] ) );
  AND2X1_RVT U400 ( .A1(n84), .A2(n48), .Y(\ab[3][15] ) );
  AND2X1_RVT U401 ( .A1(n84), .A2(n45), .Y(\ab[3][14] ) );
  AND2X1_RVT U402 ( .A1(n84), .A2(n42), .Y(\ab[3][13] ) );
  AND2X1_RVT U403 ( .A1(n84), .A2(n39), .Y(\ab[3][12] ) );
  AND2X1_RVT U404 ( .A1(n84), .A2(n36), .Y(\ab[3][11] ) );
  AND2X1_RVT U405 ( .A1(n84), .A2(n33), .Y(\ab[3][10] ) );
  AND2X1_RVT U406 ( .A1(n84), .A2(n3), .Y(\ab[3][0] ) );
  AND2X1_RVT U407 ( .A1(n82), .A2(n30), .Y(\ab[2][9] ) );
  AND2X1_RVT U408 ( .A1(n82), .A2(n27), .Y(\ab[2][8] ) );
  AND2X1_RVT U409 ( .A1(n82), .A2(n24), .Y(\ab[2][7] ) );
  AND2X1_RVT U410 ( .A1(n82), .A2(n21), .Y(\ab[2][6] ) );
  AND2X1_RVT U411 ( .A1(n82), .A2(n18), .Y(\ab[2][5] ) );
  AND2X1_RVT U412 ( .A1(n82), .A2(n15), .Y(\ab[2][4] ) );
  AND2X1_RVT U413 ( .A1(n82), .A2(n12), .Y(\ab[2][3] ) );
  AND2X1_RVT U414 ( .A1(n82), .A2(n9), .Y(\ab[2][2] ) );
  AND2X1_RVT U415 ( .A1(n82), .A2(n72), .Y(\ab[2][23] ) );
  AND2X1_RVT U416 ( .A1(n82), .A2(n69), .Y(\ab[2][22] ) );
  AND2X1_RVT U417 ( .A1(n82), .A2(n66), .Y(\ab[2][21] ) );
  AND2X1_RVT U418 ( .A1(n82), .A2(n63), .Y(\ab[2][20] ) );
  AND2X1_RVT U419 ( .A1(n81), .A2(n6), .Y(\ab[2][1] ) );
  AND2X1_RVT U420 ( .A1(n81), .A2(n60), .Y(\ab[2][19] ) );
  AND2X1_RVT U421 ( .A1(n81), .A2(n57), .Y(\ab[2][18] ) );
  AND2X1_RVT U422 ( .A1(n81), .A2(n54), .Y(\ab[2][17] ) );
  AND2X1_RVT U423 ( .A1(n81), .A2(n51), .Y(\ab[2][16] ) );
  AND2X1_RVT U424 ( .A1(n81), .A2(n48), .Y(\ab[2][15] ) );
  AND2X1_RVT U425 ( .A1(n81), .A2(n45), .Y(\ab[2][14] ) );
  AND2X1_RVT U426 ( .A1(n81), .A2(n42), .Y(\ab[2][13] ) );
  AND2X1_RVT U427 ( .A1(n81), .A2(n39), .Y(\ab[2][12] ) );
  AND2X1_RVT U428 ( .A1(n81), .A2(n36), .Y(\ab[2][11] ) );
  AND2X1_RVT U429 ( .A1(n81), .A2(n33), .Y(\ab[2][10] ) );
  AND2X1_RVT U430 ( .A1(n81), .A2(n3), .Y(\ab[2][0] ) );
  AND2X1_RVT U431 ( .A1(n145), .A2(n30), .Y(\ab[23][9] ) );
  AND2X1_RVT U432 ( .A1(n145), .A2(n27), .Y(\ab[23][8] ) );
  AND2X1_RVT U433 ( .A1(n145), .A2(n24), .Y(\ab[23][7] ) );
  AND2X1_RVT U434 ( .A1(n145), .A2(n21), .Y(\ab[23][6] ) );
  AND2X1_RVT U435 ( .A1(n145), .A2(n18), .Y(\ab[23][5] ) );
  AND2X1_RVT U436 ( .A1(n145), .A2(n15), .Y(\ab[23][4] ) );
  AND2X1_RVT U437 ( .A1(n145), .A2(n12), .Y(\ab[23][3] ) );
  AND2X1_RVT U438 ( .A1(n145), .A2(n9), .Y(\ab[23][2] ) );
  AND2X1_RVT U439 ( .A1(n145), .A2(n72), .Y(\ab[23][23] ) );
  AND2X1_RVT U440 ( .A1(n145), .A2(n69), .Y(\ab[23][22] ) );
  AND2X1_RVT U441 ( .A1(n145), .A2(n66), .Y(\ab[23][21] ) );
  AND2X1_RVT U442 ( .A1(n145), .A2(n63), .Y(\ab[23][20] ) );
  AND2X1_RVT U443 ( .A1(n144), .A2(n6), .Y(\ab[23][1] ) );
  AND2X1_RVT U444 ( .A1(n144), .A2(n60), .Y(\ab[23][19] ) );
  AND2X1_RVT U445 ( .A1(n144), .A2(n57), .Y(\ab[23][18] ) );
  AND2X1_RVT U446 ( .A1(n144), .A2(n54), .Y(\ab[23][17] ) );
  AND2X1_RVT U447 ( .A1(n144), .A2(n51), .Y(\ab[23][16] ) );
  AND2X1_RVT U448 ( .A1(n144), .A2(n48), .Y(\ab[23][15] ) );
  AND2X1_RVT U449 ( .A1(n144), .A2(n45), .Y(\ab[23][14] ) );
  AND2X1_RVT U450 ( .A1(n144), .A2(n42), .Y(\ab[23][13] ) );
  AND2X1_RVT U451 ( .A1(n144), .A2(n39), .Y(\ab[23][12] ) );
  AND2X1_RVT U452 ( .A1(n144), .A2(n36), .Y(\ab[23][11] ) );
  AND2X1_RVT U453 ( .A1(n144), .A2(n33), .Y(\ab[23][10] ) );
  AND2X1_RVT U454 ( .A1(n144), .A2(n3), .Y(\ab[23][0] ) );
  AND2X1_RVT U455 ( .A1(n142), .A2(n30), .Y(\ab[22][9] ) );
  AND2X1_RVT U456 ( .A1(n142), .A2(n27), .Y(\ab[22][8] ) );
  AND2X1_RVT U457 ( .A1(n142), .A2(n24), .Y(\ab[22][7] ) );
  AND2X1_RVT U458 ( .A1(n142), .A2(n21), .Y(\ab[22][6] ) );
  AND2X1_RVT U459 ( .A1(n142), .A2(n18), .Y(\ab[22][5] ) );
  AND2X1_RVT U460 ( .A1(n142), .A2(n15), .Y(\ab[22][4] ) );
  AND2X1_RVT U461 ( .A1(n142), .A2(n12), .Y(\ab[22][3] ) );
  AND2X1_RVT U462 ( .A1(n142), .A2(n9), .Y(\ab[22][2] ) );
  AND2X1_RVT U463 ( .A1(n142), .A2(n72), .Y(\ab[22][23] ) );
  AND2X1_RVT U464 ( .A1(n142), .A2(n69), .Y(\ab[22][22] ) );
  AND2X1_RVT U465 ( .A1(n142), .A2(n66), .Y(\ab[22][21] ) );
  AND2X1_RVT U466 ( .A1(n142), .A2(n63), .Y(\ab[22][20] ) );
  AND2X1_RVT U467 ( .A1(n141), .A2(n6), .Y(\ab[22][1] ) );
  AND2X1_RVT U468 ( .A1(n141), .A2(n60), .Y(\ab[22][19] ) );
  AND2X1_RVT U469 ( .A1(n141), .A2(n57), .Y(\ab[22][18] ) );
  AND2X1_RVT U470 ( .A1(n141), .A2(n54), .Y(\ab[22][17] ) );
  AND2X1_RVT U471 ( .A1(n141), .A2(n51), .Y(\ab[22][16] ) );
  AND2X1_RVT U472 ( .A1(n141), .A2(n48), .Y(\ab[22][15] ) );
  AND2X1_RVT U473 ( .A1(n141), .A2(n45), .Y(\ab[22][14] ) );
  AND2X1_RVT U474 ( .A1(n141), .A2(n42), .Y(\ab[22][13] ) );
  AND2X1_RVT U475 ( .A1(n141), .A2(n39), .Y(\ab[22][12] ) );
  AND2X1_RVT U476 ( .A1(n141), .A2(n36), .Y(\ab[22][11] ) );
  AND2X1_RVT U477 ( .A1(n141), .A2(n33), .Y(\ab[22][10] ) );
  AND2X1_RVT U478 ( .A1(n141), .A2(n3), .Y(\ab[22][0] ) );
  AND2X1_RVT U479 ( .A1(n139), .A2(n30), .Y(\ab[21][9] ) );
  AND2X1_RVT U480 ( .A1(n139), .A2(n27), .Y(\ab[21][8] ) );
  AND2X1_RVT U481 ( .A1(n139), .A2(n24), .Y(\ab[21][7] ) );
  AND2X1_RVT U482 ( .A1(n139), .A2(n21), .Y(\ab[21][6] ) );
  AND2X1_RVT U483 ( .A1(n139), .A2(n18), .Y(\ab[21][5] ) );
  AND2X1_RVT U484 ( .A1(n139), .A2(n15), .Y(\ab[21][4] ) );
  AND2X1_RVT U485 ( .A1(n139), .A2(n12), .Y(\ab[21][3] ) );
  AND2X1_RVT U486 ( .A1(n139), .A2(n9), .Y(\ab[21][2] ) );
  AND2X1_RVT U487 ( .A1(n139), .A2(n72), .Y(\ab[21][23] ) );
  AND2X1_RVT U488 ( .A1(n139), .A2(n69), .Y(\ab[21][22] ) );
  AND2X1_RVT U489 ( .A1(n139), .A2(n66), .Y(\ab[21][21] ) );
  AND2X1_RVT U490 ( .A1(n139), .A2(n63), .Y(\ab[21][20] ) );
  AND2X1_RVT U491 ( .A1(n138), .A2(n6), .Y(\ab[21][1] ) );
  AND2X1_RVT U492 ( .A1(n138), .A2(n60), .Y(\ab[21][19] ) );
  AND2X1_RVT U493 ( .A1(n138), .A2(n57), .Y(\ab[21][18] ) );
  AND2X1_RVT U494 ( .A1(n138), .A2(n54), .Y(\ab[21][17] ) );
  AND2X1_RVT U495 ( .A1(n138), .A2(n51), .Y(\ab[21][16] ) );
  AND2X1_RVT U496 ( .A1(n138), .A2(n48), .Y(\ab[21][15] ) );
  AND2X1_RVT U497 ( .A1(n138), .A2(n45), .Y(\ab[21][14] ) );
  AND2X1_RVT U498 ( .A1(n138), .A2(n42), .Y(\ab[21][13] ) );
  AND2X1_RVT U499 ( .A1(n138), .A2(n39), .Y(\ab[21][12] ) );
  AND2X1_RVT U500 ( .A1(n138), .A2(n36), .Y(\ab[21][11] ) );
  AND2X1_RVT U501 ( .A1(n138), .A2(n33), .Y(\ab[21][10] ) );
  AND2X1_RVT U502 ( .A1(n138), .A2(n3), .Y(\ab[21][0] ) );
  AND2X1_RVT U503 ( .A1(n136), .A2(n30), .Y(\ab[20][9] ) );
  AND2X1_RVT U504 ( .A1(n136), .A2(n27), .Y(\ab[20][8] ) );
  AND2X1_RVT U505 ( .A1(n136), .A2(n24), .Y(\ab[20][7] ) );
  AND2X1_RVT U506 ( .A1(n136), .A2(n21), .Y(\ab[20][6] ) );
  AND2X1_RVT U507 ( .A1(n136), .A2(n18), .Y(\ab[20][5] ) );
  AND2X1_RVT U508 ( .A1(n136), .A2(n15), .Y(\ab[20][4] ) );
  AND2X1_RVT U509 ( .A1(n136), .A2(n12), .Y(\ab[20][3] ) );
  AND2X1_RVT U510 ( .A1(n136), .A2(n9), .Y(\ab[20][2] ) );
  AND2X1_RVT U511 ( .A1(n136), .A2(n72), .Y(\ab[20][23] ) );
  AND2X1_RVT U512 ( .A1(n136), .A2(n69), .Y(\ab[20][22] ) );
  AND2X1_RVT U513 ( .A1(n136), .A2(n66), .Y(\ab[20][21] ) );
  AND2X1_RVT U514 ( .A1(n136), .A2(n63), .Y(\ab[20][20] ) );
  AND2X1_RVT U515 ( .A1(n135), .A2(n6), .Y(\ab[20][1] ) );
  AND2X1_RVT U516 ( .A1(n135), .A2(n60), .Y(\ab[20][19] ) );
  AND2X1_RVT U517 ( .A1(n135), .A2(n57), .Y(\ab[20][18] ) );
  AND2X1_RVT U518 ( .A1(n135), .A2(n54), .Y(\ab[20][17] ) );
  AND2X1_RVT U519 ( .A1(n135), .A2(n51), .Y(\ab[20][16] ) );
  AND2X1_RVT U520 ( .A1(n135), .A2(n48), .Y(\ab[20][15] ) );
  AND2X1_RVT U521 ( .A1(n135), .A2(n45), .Y(\ab[20][14] ) );
  AND2X1_RVT U522 ( .A1(n135), .A2(n42), .Y(\ab[20][13] ) );
  AND2X1_RVT U523 ( .A1(n135), .A2(n39), .Y(\ab[20][12] ) );
  AND2X1_RVT U524 ( .A1(n135), .A2(n36), .Y(\ab[20][11] ) );
  AND2X1_RVT U525 ( .A1(n135), .A2(n33), .Y(\ab[20][10] ) );
  AND2X1_RVT U526 ( .A1(n135), .A2(n3), .Y(\ab[20][0] ) );
  AND2X1_RVT U527 ( .A1(n79), .A2(n30), .Y(\ab[1][9] ) );
  AND2X1_RVT U528 ( .A1(n79), .A2(n27), .Y(\ab[1][8] ) );
  AND2X1_RVT U529 ( .A1(n79), .A2(n24), .Y(\ab[1][7] ) );
  AND2X1_RVT U530 ( .A1(n79), .A2(n21), .Y(\ab[1][6] ) );
  AND2X1_RVT U531 ( .A1(n79), .A2(n18), .Y(\ab[1][5] ) );
  AND2X1_RVT U532 ( .A1(n79), .A2(n15), .Y(\ab[1][4] ) );
  AND2X1_RVT U533 ( .A1(n79), .A2(n12), .Y(\ab[1][3] ) );
  AND2X1_RVT U534 ( .A1(n79), .A2(n9), .Y(\ab[1][2] ) );
  AND2X1_RVT U535 ( .A1(n79), .A2(n72), .Y(\ab[1][23] ) );
  AND2X1_RVT U536 ( .A1(n79), .A2(n69), .Y(\ab[1][22] ) );
  AND2X1_RVT U537 ( .A1(n79), .A2(n66), .Y(\ab[1][21] ) );
  AND2X1_RVT U538 ( .A1(n79), .A2(n63), .Y(\ab[1][20] ) );
  AND2X1_RVT U539 ( .A1(n78), .A2(n6), .Y(\ab[1][1] ) );
  AND2X1_RVT U540 ( .A1(n78), .A2(n60), .Y(\ab[1][19] ) );
  AND2X1_RVT U541 ( .A1(n78), .A2(n57), .Y(\ab[1][18] ) );
  AND2X1_RVT U542 ( .A1(n78), .A2(n54), .Y(\ab[1][17] ) );
  AND2X1_RVT U543 ( .A1(n78), .A2(n51), .Y(\ab[1][16] ) );
  AND2X1_RVT U544 ( .A1(n78), .A2(n48), .Y(\ab[1][15] ) );
  AND2X1_RVT U545 ( .A1(n78), .A2(n45), .Y(\ab[1][14] ) );
  AND2X1_RVT U546 ( .A1(n78), .A2(n42), .Y(\ab[1][13] ) );
  AND2X1_RVT U547 ( .A1(n78), .A2(n39), .Y(\ab[1][12] ) );
  AND2X1_RVT U548 ( .A1(n78), .A2(n36), .Y(\ab[1][11] ) );
  AND2X1_RVT U549 ( .A1(n78), .A2(n33), .Y(\ab[1][10] ) );
  AND2X1_RVT U550 ( .A1(n78), .A2(n3), .Y(\ab[1][0] ) );
  AND2X1_RVT U551 ( .A1(n133), .A2(n30), .Y(\ab[19][9] ) );
  AND2X1_RVT U552 ( .A1(n133), .A2(n27), .Y(\ab[19][8] ) );
  AND2X1_RVT U553 ( .A1(n133), .A2(n24), .Y(\ab[19][7] ) );
  AND2X1_RVT U554 ( .A1(n133), .A2(n21), .Y(\ab[19][6] ) );
  AND2X1_RVT U555 ( .A1(n133), .A2(n18), .Y(\ab[19][5] ) );
  AND2X1_RVT U556 ( .A1(n133), .A2(n15), .Y(\ab[19][4] ) );
  AND2X1_RVT U557 ( .A1(n133), .A2(n12), .Y(\ab[19][3] ) );
  AND2X1_RVT U558 ( .A1(n133), .A2(n9), .Y(\ab[19][2] ) );
  AND2X1_RVT U559 ( .A1(n133), .A2(n72), .Y(\ab[19][23] ) );
  AND2X1_RVT U560 ( .A1(n133), .A2(n69), .Y(\ab[19][22] ) );
  AND2X1_RVT U561 ( .A1(n133), .A2(n66), .Y(\ab[19][21] ) );
  AND2X1_RVT U562 ( .A1(n133), .A2(n63), .Y(\ab[19][20] ) );
  AND2X1_RVT U563 ( .A1(n132), .A2(n6), .Y(\ab[19][1] ) );
  AND2X1_RVT U564 ( .A1(n132), .A2(n60), .Y(\ab[19][19] ) );
  AND2X1_RVT U565 ( .A1(n132), .A2(n57), .Y(\ab[19][18] ) );
  AND2X1_RVT U566 ( .A1(n132), .A2(n54), .Y(\ab[19][17] ) );
  AND2X1_RVT U567 ( .A1(n132), .A2(n51), .Y(\ab[19][16] ) );
  AND2X1_RVT U568 ( .A1(n132), .A2(n48), .Y(\ab[19][15] ) );
  AND2X1_RVT U569 ( .A1(n132), .A2(n45), .Y(\ab[19][14] ) );
  AND2X1_RVT U570 ( .A1(n132), .A2(n42), .Y(\ab[19][13] ) );
  AND2X1_RVT U571 ( .A1(n132), .A2(n39), .Y(\ab[19][12] ) );
  AND2X1_RVT U572 ( .A1(n132), .A2(n36), .Y(\ab[19][11] ) );
  AND2X1_RVT U573 ( .A1(n132), .A2(n33), .Y(\ab[19][10] ) );
  AND2X1_RVT U574 ( .A1(n132), .A2(n3), .Y(\ab[19][0] ) );
  AND2X1_RVT U575 ( .A1(n130), .A2(n31), .Y(\ab[18][9] ) );
  AND2X1_RVT U576 ( .A1(n130), .A2(n28), .Y(\ab[18][8] ) );
  AND2X1_RVT U577 ( .A1(n130), .A2(n25), .Y(\ab[18][7] ) );
  AND2X1_RVT U578 ( .A1(n130), .A2(n22), .Y(\ab[18][6] ) );
  AND2X1_RVT U579 ( .A1(n130), .A2(n19), .Y(\ab[18][5] ) );
  AND2X1_RVT U580 ( .A1(n130), .A2(n16), .Y(\ab[18][4] ) );
  AND2X1_RVT U581 ( .A1(n130), .A2(n13), .Y(\ab[18][3] ) );
  AND2X1_RVT U582 ( .A1(n130), .A2(n10), .Y(\ab[18][2] ) );
  AND2X1_RVT U583 ( .A1(n130), .A2(n73), .Y(\ab[18][23] ) );
  AND2X1_RVT U584 ( .A1(n130), .A2(n70), .Y(\ab[18][22] ) );
  AND2X1_RVT U585 ( .A1(n130), .A2(n67), .Y(\ab[18][21] ) );
  AND2X1_RVT U586 ( .A1(n130), .A2(n64), .Y(\ab[18][20] ) );
  AND2X1_RVT U587 ( .A1(n129), .A2(n7), .Y(\ab[18][1] ) );
  AND2X1_RVT U588 ( .A1(n129), .A2(n61), .Y(\ab[18][19] ) );
  AND2X1_RVT U589 ( .A1(n129), .A2(n58), .Y(\ab[18][18] ) );
  AND2X1_RVT U590 ( .A1(n129), .A2(n55), .Y(\ab[18][17] ) );
  AND2X1_RVT U591 ( .A1(n129), .A2(n52), .Y(\ab[18][16] ) );
  AND2X1_RVT U592 ( .A1(n129), .A2(n49), .Y(\ab[18][15] ) );
  AND2X1_RVT U593 ( .A1(n129), .A2(n46), .Y(\ab[18][14] ) );
  AND2X1_RVT U594 ( .A1(n129), .A2(n43), .Y(\ab[18][13] ) );
  AND2X1_RVT U595 ( .A1(n129), .A2(n40), .Y(\ab[18][12] ) );
  AND2X1_RVT U596 ( .A1(n129), .A2(n37), .Y(\ab[18][11] ) );
  AND2X1_RVT U597 ( .A1(n129), .A2(n34), .Y(\ab[18][10] ) );
  AND2X1_RVT U598 ( .A1(n129), .A2(n4), .Y(\ab[18][0] ) );
  AND2X1_RVT U599 ( .A1(n127), .A2(n31), .Y(\ab[17][9] ) );
  AND2X1_RVT U600 ( .A1(n127), .A2(n28), .Y(\ab[17][8] ) );
  AND2X1_RVT U601 ( .A1(n127), .A2(n25), .Y(\ab[17][7] ) );
  AND2X1_RVT U602 ( .A1(n127), .A2(n22), .Y(\ab[17][6] ) );
  AND2X1_RVT U603 ( .A1(n127), .A2(n19), .Y(\ab[17][5] ) );
  AND2X1_RVT U604 ( .A1(n127), .A2(n16), .Y(\ab[17][4] ) );
  AND2X1_RVT U605 ( .A1(n127), .A2(n13), .Y(\ab[17][3] ) );
  AND2X1_RVT U606 ( .A1(n127), .A2(n10), .Y(\ab[17][2] ) );
  AND2X1_RVT U607 ( .A1(n127), .A2(n73), .Y(\ab[17][23] ) );
  AND2X1_RVT U608 ( .A1(n127), .A2(n70), .Y(\ab[17][22] ) );
  AND2X1_RVT U609 ( .A1(n127), .A2(n67), .Y(\ab[17][21] ) );
  AND2X1_RVT U610 ( .A1(n127), .A2(n64), .Y(\ab[17][20] ) );
  AND2X1_RVT U611 ( .A1(n126), .A2(n7), .Y(\ab[17][1] ) );
  AND2X1_RVT U612 ( .A1(n126), .A2(n61), .Y(\ab[17][19] ) );
  AND2X1_RVT U613 ( .A1(n126), .A2(n58), .Y(\ab[17][18] ) );
  AND2X1_RVT U614 ( .A1(n126), .A2(n55), .Y(\ab[17][17] ) );
  AND2X1_RVT U615 ( .A1(n126), .A2(n52), .Y(\ab[17][16] ) );
  AND2X1_RVT U616 ( .A1(n126), .A2(n49), .Y(\ab[17][15] ) );
  AND2X1_RVT U617 ( .A1(n126), .A2(n46), .Y(\ab[17][14] ) );
  AND2X1_RVT U618 ( .A1(n126), .A2(n43), .Y(\ab[17][13] ) );
  AND2X1_RVT U619 ( .A1(n126), .A2(n40), .Y(\ab[17][12] ) );
  AND2X1_RVT U620 ( .A1(n126), .A2(n37), .Y(\ab[17][11] ) );
  AND2X1_RVT U621 ( .A1(n126), .A2(n34), .Y(\ab[17][10] ) );
  AND2X1_RVT U622 ( .A1(n126), .A2(n4), .Y(\ab[17][0] ) );
  AND2X1_RVT U623 ( .A1(n124), .A2(n31), .Y(\ab[16][9] ) );
  AND2X1_RVT U624 ( .A1(n124), .A2(n28), .Y(\ab[16][8] ) );
  AND2X1_RVT U625 ( .A1(n124), .A2(n25), .Y(\ab[16][7] ) );
  AND2X1_RVT U626 ( .A1(n124), .A2(n22), .Y(\ab[16][6] ) );
  AND2X1_RVT U627 ( .A1(n124), .A2(n19), .Y(\ab[16][5] ) );
  AND2X1_RVT U628 ( .A1(n124), .A2(n16), .Y(\ab[16][4] ) );
  AND2X1_RVT U629 ( .A1(n124), .A2(n13), .Y(\ab[16][3] ) );
  AND2X1_RVT U630 ( .A1(n124), .A2(n10), .Y(\ab[16][2] ) );
  AND2X1_RVT U631 ( .A1(n124), .A2(n73), .Y(\ab[16][23] ) );
  AND2X1_RVT U632 ( .A1(n124), .A2(n70), .Y(\ab[16][22] ) );
  AND2X1_RVT U633 ( .A1(n124), .A2(n67), .Y(\ab[16][21] ) );
  AND2X1_RVT U634 ( .A1(n124), .A2(n64), .Y(\ab[16][20] ) );
  AND2X1_RVT U635 ( .A1(n123), .A2(n7), .Y(\ab[16][1] ) );
  AND2X1_RVT U636 ( .A1(n123), .A2(n61), .Y(\ab[16][19] ) );
  AND2X1_RVT U637 ( .A1(n123), .A2(n58), .Y(\ab[16][18] ) );
  AND2X1_RVT U638 ( .A1(n123), .A2(n55), .Y(\ab[16][17] ) );
  AND2X1_RVT U639 ( .A1(n123), .A2(n52), .Y(\ab[16][16] ) );
  AND2X1_RVT U640 ( .A1(n123), .A2(n49), .Y(\ab[16][15] ) );
  AND2X1_RVT U641 ( .A1(n123), .A2(n46), .Y(\ab[16][14] ) );
  AND2X1_RVT U642 ( .A1(n123), .A2(n43), .Y(\ab[16][13] ) );
  AND2X1_RVT U643 ( .A1(n123), .A2(n40), .Y(\ab[16][12] ) );
  AND2X1_RVT U644 ( .A1(n123), .A2(n37), .Y(\ab[16][11] ) );
  AND2X1_RVT U645 ( .A1(n123), .A2(n34), .Y(\ab[16][10] ) );
  AND2X1_RVT U646 ( .A1(n123), .A2(n4), .Y(\ab[16][0] ) );
  AND2X1_RVT U647 ( .A1(n121), .A2(n31), .Y(\ab[15][9] ) );
  AND2X1_RVT U648 ( .A1(n121), .A2(n28), .Y(\ab[15][8] ) );
  AND2X1_RVT U649 ( .A1(n121), .A2(n25), .Y(\ab[15][7] ) );
  AND2X1_RVT U650 ( .A1(n121), .A2(n22), .Y(\ab[15][6] ) );
  AND2X1_RVT U651 ( .A1(n121), .A2(n19), .Y(\ab[15][5] ) );
  AND2X1_RVT U652 ( .A1(n121), .A2(n16), .Y(\ab[15][4] ) );
  AND2X1_RVT U653 ( .A1(n121), .A2(n13), .Y(\ab[15][3] ) );
  AND2X1_RVT U654 ( .A1(n121), .A2(n10), .Y(\ab[15][2] ) );
  AND2X1_RVT U655 ( .A1(n121), .A2(n73), .Y(\ab[15][23] ) );
  AND2X1_RVT U656 ( .A1(n121), .A2(n70), .Y(\ab[15][22] ) );
  AND2X1_RVT U657 ( .A1(n121), .A2(n67), .Y(\ab[15][21] ) );
  AND2X1_RVT U658 ( .A1(n121), .A2(n64), .Y(\ab[15][20] ) );
  AND2X1_RVT U659 ( .A1(n120), .A2(n7), .Y(\ab[15][1] ) );
  AND2X1_RVT U660 ( .A1(n120), .A2(n61), .Y(\ab[15][19] ) );
  AND2X1_RVT U661 ( .A1(n120), .A2(n58), .Y(\ab[15][18] ) );
  AND2X1_RVT U662 ( .A1(n120), .A2(n55), .Y(\ab[15][17] ) );
  AND2X1_RVT U663 ( .A1(n120), .A2(n52), .Y(\ab[15][16] ) );
  AND2X1_RVT U664 ( .A1(n120), .A2(n49), .Y(\ab[15][15] ) );
  AND2X1_RVT U665 ( .A1(n120), .A2(n46), .Y(\ab[15][14] ) );
  AND2X1_RVT U666 ( .A1(n120), .A2(n43), .Y(\ab[15][13] ) );
  AND2X1_RVT U667 ( .A1(n120), .A2(n40), .Y(\ab[15][12] ) );
  AND2X1_RVT U668 ( .A1(n120), .A2(n37), .Y(\ab[15][11] ) );
  AND2X1_RVT U669 ( .A1(n120), .A2(n34), .Y(\ab[15][10] ) );
  AND2X1_RVT U670 ( .A1(n120), .A2(n4), .Y(\ab[15][0] ) );
  AND2X1_RVT U671 ( .A1(n118), .A2(n31), .Y(\ab[14][9] ) );
  AND2X1_RVT U672 ( .A1(n118), .A2(n28), .Y(\ab[14][8] ) );
  AND2X1_RVT U673 ( .A1(n118), .A2(n25), .Y(\ab[14][7] ) );
  AND2X1_RVT U674 ( .A1(n118), .A2(n22), .Y(\ab[14][6] ) );
  AND2X1_RVT U675 ( .A1(n118), .A2(n19), .Y(\ab[14][5] ) );
  AND2X1_RVT U676 ( .A1(n118), .A2(n16), .Y(\ab[14][4] ) );
  AND2X1_RVT U677 ( .A1(n118), .A2(n13), .Y(\ab[14][3] ) );
  AND2X1_RVT U678 ( .A1(n118), .A2(n10), .Y(\ab[14][2] ) );
  AND2X1_RVT U679 ( .A1(n118), .A2(n73), .Y(\ab[14][23] ) );
  AND2X1_RVT U680 ( .A1(n118), .A2(n70), .Y(\ab[14][22] ) );
  AND2X1_RVT U681 ( .A1(n118), .A2(n67), .Y(\ab[14][21] ) );
  AND2X1_RVT U682 ( .A1(n118), .A2(n64), .Y(\ab[14][20] ) );
  AND2X1_RVT U683 ( .A1(n117), .A2(n7), .Y(\ab[14][1] ) );
  AND2X1_RVT U684 ( .A1(n117), .A2(n61), .Y(\ab[14][19] ) );
  AND2X1_RVT U685 ( .A1(n117), .A2(n58), .Y(\ab[14][18] ) );
  AND2X1_RVT U686 ( .A1(n117), .A2(n55), .Y(\ab[14][17] ) );
  AND2X1_RVT U687 ( .A1(n117), .A2(n52), .Y(\ab[14][16] ) );
  AND2X1_RVT U688 ( .A1(n117), .A2(n49), .Y(\ab[14][15] ) );
  AND2X1_RVT U689 ( .A1(n117), .A2(n46), .Y(\ab[14][14] ) );
  AND2X1_RVT U690 ( .A1(n117), .A2(n43), .Y(\ab[14][13] ) );
  AND2X1_RVT U691 ( .A1(n117), .A2(n40), .Y(\ab[14][12] ) );
  AND2X1_RVT U692 ( .A1(n117), .A2(n37), .Y(\ab[14][11] ) );
  AND2X1_RVT U693 ( .A1(n117), .A2(n34), .Y(\ab[14][10] ) );
  AND2X1_RVT U694 ( .A1(n117), .A2(n4), .Y(\ab[14][0] ) );
  AND2X1_RVT U695 ( .A1(n115), .A2(n31), .Y(\ab[13][9] ) );
  AND2X1_RVT U696 ( .A1(n115), .A2(n28), .Y(\ab[13][8] ) );
  AND2X1_RVT U697 ( .A1(n115), .A2(n25), .Y(\ab[13][7] ) );
  AND2X1_RVT U698 ( .A1(n115), .A2(n22), .Y(\ab[13][6] ) );
  AND2X1_RVT U699 ( .A1(n115), .A2(n19), .Y(\ab[13][5] ) );
  AND2X1_RVT U700 ( .A1(n115), .A2(n16), .Y(\ab[13][4] ) );
  AND2X1_RVT U701 ( .A1(n115), .A2(n13), .Y(\ab[13][3] ) );
  AND2X1_RVT U702 ( .A1(n115), .A2(n10), .Y(\ab[13][2] ) );
  AND2X1_RVT U703 ( .A1(n115), .A2(n73), .Y(\ab[13][23] ) );
  AND2X1_RVT U704 ( .A1(n115), .A2(n70), .Y(\ab[13][22] ) );
  AND2X1_RVT U705 ( .A1(n115), .A2(n67), .Y(\ab[13][21] ) );
  AND2X1_RVT U706 ( .A1(n115), .A2(n64), .Y(\ab[13][20] ) );
  AND2X1_RVT U707 ( .A1(n114), .A2(n7), .Y(\ab[13][1] ) );
  AND2X1_RVT U708 ( .A1(n114), .A2(n61), .Y(\ab[13][19] ) );
  AND2X1_RVT U709 ( .A1(n114), .A2(n58), .Y(\ab[13][18] ) );
  AND2X1_RVT U710 ( .A1(n114), .A2(n55), .Y(\ab[13][17] ) );
  AND2X1_RVT U711 ( .A1(n114), .A2(n52), .Y(\ab[13][16] ) );
  AND2X1_RVT U712 ( .A1(n114), .A2(n49), .Y(\ab[13][15] ) );
  AND2X1_RVT U713 ( .A1(n114), .A2(n46), .Y(\ab[13][14] ) );
  AND2X1_RVT U714 ( .A1(n114), .A2(n43), .Y(\ab[13][13] ) );
  AND2X1_RVT U715 ( .A1(n114), .A2(n40), .Y(\ab[13][12] ) );
  AND2X1_RVT U716 ( .A1(n114), .A2(n37), .Y(\ab[13][11] ) );
  AND2X1_RVT U717 ( .A1(n114), .A2(n34), .Y(\ab[13][10] ) );
  AND2X1_RVT U718 ( .A1(n114), .A2(n4), .Y(\ab[13][0] ) );
  AND2X1_RVT U719 ( .A1(n112), .A2(n31), .Y(\ab[12][9] ) );
  AND2X1_RVT U720 ( .A1(n112), .A2(n28), .Y(\ab[12][8] ) );
  AND2X1_RVT U721 ( .A1(n112), .A2(n25), .Y(\ab[12][7] ) );
  AND2X1_RVT U722 ( .A1(n112), .A2(n22), .Y(\ab[12][6] ) );
  AND2X1_RVT U723 ( .A1(n112), .A2(n19), .Y(\ab[12][5] ) );
  AND2X1_RVT U724 ( .A1(n112), .A2(n16), .Y(\ab[12][4] ) );
  AND2X1_RVT U725 ( .A1(n112), .A2(n13), .Y(\ab[12][3] ) );
  AND2X1_RVT U726 ( .A1(n112), .A2(n10), .Y(\ab[12][2] ) );
  AND2X1_RVT U727 ( .A1(n112), .A2(n73), .Y(\ab[12][23] ) );
  AND2X1_RVT U728 ( .A1(n112), .A2(n70), .Y(\ab[12][22] ) );
  AND2X1_RVT U729 ( .A1(n112), .A2(n67), .Y(\ab[12][21] ) );
  AND2X1_RVT U730 ( .A1(n112), .A2(n64), .Y(\ab[12][20] ) );
  AND2X1_RVT U731 ( .A1(n111), .A2(n7), .Y(\ab[12][1] ) );
  AND2X1_RVT U732 ( .A1(n111), .A2(n61), .Y(\ab[12][19] ) );
  AND2X1_RVT U733 ( .A1(n111), .A2(n58), .Y(\ab[12][18] ) );
  AND2X1_RVT U734 ( .A1(n111), .A2(n55), .Y(\ab[12][17] ) );
  AND2X1_RVT U735 ( .A1(n111), .A2(n52), .Y(\ab[12][16] ) );
  AND2X1_RVT U736 ( .A1(n111), .A2(n49), .Y(\ab[12][15] ) );
  AND2X1_RVT U737 ( .A1(n111), .A2(n46), .Y(\ab[12][14] ) );
  AND2X1_RVT U738 ( .A1(n111), .A2(n43), .Y(\ab[12][13] ) );
  AND2X1_RVT U739 ( .A1(n111), .A2(n40), .Y(\ab[12][12] ) );
  AND2X1_RVT U740 ( .A1(n111), .A2(n37), .Y(\ab[12][11] ) );
  AND2X1_RVT U741 ( .A1(n111), .A2(n34), .Y(\ab[12][10] ) );
  AND2X1_RVT U742 ( .A1(n111), .A2(n4), .Y(\ab[12][0] ) );
  AND2X1_RVT U743 ( .A1(n109), .A2(n31), .Y(\ab[11][9] ) );
  AND2X1_RVT U744 ( .A1(n109), .A2(n28), .Y(\ab[11][8] ) );
  AND2X1_RVT U745 ( .A1(n109), .A2(n25), .Y(\ab[11][7] ) );
  AND2X1_RVT U746 ( .A1(n109), .A2(n22), .Y(\ab[11][6] ) );
  AND2X1_RVT U747 ( .A1(n109), .A2(n19), .Y(\ab[11][5] ) );
  AND2X1_RVT U748 ( .A1(n109), .A2(n16), .Y(\ab[11][4] ) );
  AND2X1_RVT U749 ( .A1(n109), .A2(n13), .Y(\ab[11][3] ) );
  AND2X1_RVT U750 ( .A1(n109), .A2(n10), .Y(\ab[11][2] ) );
  AND2X1_RVT U751 ( .A1(n109), .A2(n73), .Y(\ab[11][23] ) );
  AND2X1_RVT U752 ( .A1(n109), .A2(n70), .Y(\ab[11][22] ) );
  AND2X1_RVT U753 ( .A1(n109), .A2(n67), .Y(\ab[11][21] ) );
  AND2X1_RVT U754 ( .A1(n109), .A2(n64), .Y(\ab[11][20] ) );
  AND2X1_RVT U755 ( .A1(n108), .A2(n7), .Y(\ab[11][1] ) );
  AND2X1_RVT U756 ( .A1(n108), .A2(n61), .Y(\ab[11][19] ) );
  AND2X1_RVT U757 ( .A1(n108), .A2(n58), .Y(\ab[11][18] ) );
  AND2X1_RVT U758 ( .A1(n108), .A2(n55), .Y(\ab[11][17] ) );
  AND2X1_RVT U759 ( .A1(n108), .A2(n52), .Y(\ab[11][16] ) );
  AND2X1_RVT U760 ( .A1(n108), .A2(n49), .Y(\ab[11][15] ) );
  AND2X1_RVT U761 ( .A1(n108), .A2(n46), .Y(\ab[11][14] ) );
  AND2X1_RVT U762 ( .A1(n108), .A2(n43), .Y(\ab[11][13] ) );
  AND2X1_RVT U763 ( .A1(n108), .A2(n40), .Y(\ab[11][12] ) );
  AND2X1_RVT U764 ( .A1(n108), .A2(n37), .Y(\ab[11][11] ) );
  AND2X1_RVT U765 ( .A1(n108), .A2(n34), .Y(\ab[11][10] ) );
  AND2X1_RVT U766 ( .A1(n108), .A2(n4), .Y(\ab[11][0] ) );
  AND2X1_RVT U767 ( .A1(n106), .A2(n31), .Y(\ab[10][9] ) );
  AND2X1_RVT U768 ( .A1(n106), .A2(n28), .Y(\ab[10][8] ) );
  AND2X1_RVT U769 ( .A1(n106), .A2(n25), .Y(\ab[10][7] ) );
  AND2X1_RVT U770 ( .A1(n106), .A2(n22), .Y(\ab[10][6] ) );
  AND2X1_RVT U771 ( .A1(n106), .A2(n19), .Y(\ab[10][5] ) );
  AND2X1_RVT U772 ( .A1(n106), .A2(n16), .Y(\ab[10][4] ) );
  AND2X1_RVT U773 ( .A1(n106), .A2(n13), .Y(\ab[10][3] ) );
  AND2X1_RVT U774 ( .A1(n106), .A2(n10), .Y(\ab[10][2] ) );
  AND2X1_RVT U775 ( .A1(n106), .A2(n73), .Y(\ab[10][23] ) );
  AND2X1_RVT U776 ( .A1(n106), .A2(n70), .Y(\ab[10][22] ) );
  AND2X1_RVT U777 ( .A1(n106), .A2(n67), .Y(\ab[10][21] ) );
  AND2X1_RVT U778 ( .A1(n106), .A2(n64), .Y(\ab[10][20] ) );
  AND2X1_RVT U779 ( .A1(n105), .A2(n7), .Y(\ab[10][1] ) );
  AND2X1_RVT U780 ( .A1(n105), .A2(n61), .Y(\ab[10][19] ) );
  AND2X1_RVT U781 ( .A1(n105), .A2(n58), .Y(\ab[10][18] ) );
  AND2X1_RVT U782 ( .A1(n105), .A2(n55), .Y(\ab[10][17] ) );
  AND2X1_RVT U783 ( .A1(n105), .A2(n52), .Y(\ab[10][16] ) );
  AND2X1_RVT U784 ( .A1(n105), .A2(n49), .Y(\ab[10][15] ) );
  AND2X1_RVT U785 ( .A1(n105), .A2(n46), .Y(\ab[10][14] ) );
  AND2X1_RVT U786 ( .A1(n105), .A2(n43), .Y(\ab[10][13] ) );
  AND2X1_RVT U787 ( .A1(n105), .A2(n40), .Y(\ab[10][12] ) );
  AND2X1_RVT U788 ( .A1(n105), .A2(n37), .Y(\ab[10][11] ) );
  AND2X1_RVT U789 ( .A1(n105), .A2(n34), .Y(\ab[10][10] ) );
  AND2X1_RVT U790 ( .A1(n105), .A2(n4), .Y(\ab[10][0] ) );
  AND2X1_RVT U791 ( .A1(n76), .A2(n31), .Y(\ab[0][9] ) );
  AND2X1_RVT U792 ( .A1(n76), .A2(n28), .Y(\ab[0][8] ) );
  AND2X1_RVT U793 ( .A1(n76), .A2(n25), .Y(\ab[0][7] ) );
  AND2X1_RVT U794 ( .A1(n76), .A2(n22), .Y(\ab[0][6] ) );
  AND2X1_RVT U795 ( .A1(n76), .A2(n19), .Y(\ab[0][5] ) );
  AND2X1_RVT U796 ( .A1(n76), .A2(n16), .Y(\ab[0][4] ) );
  AND2X1_RVT U797 ( .A1(n76), .A2(n13), .Y(\ab[0][3] ) );
  AND2X1_RVT U798 ( .A1(n76), .A2(n10), .Y(\ab[0][2] ) );
  AND2X1_RVT U799 ( .A1(n76), .A2(n73), .Y(\ab[0][23] ) );
  AND2X1_RVT U800 ( .A1(n76), .A2(n70), .Y(\ab[0][22] ) );
  AND2X1_RVT U801 ( .A1(n76), .A2(n67), .Y(\ab[0][21] ) );
  AND2X1_RVT U802 ( .A1(n76), .A2(n64), .Y(\ab[0][20] ) );
  AND2X1_RVT U803 ( .A1(n75), .A2(n7), .Y(\ab[0][1] ) );
  AND2X1_RVT U804 ( .A1(n75), .A2(n61), .Y(\ab[0][19] ) );
  AND2X1_RVT U805 ( .A1(n75), .A2(n58), .Y(\ab[0][18] ) );
  AND2X1_RVT U806 ( .A1(n75), .A2(n55), .Y(\ab[0][17] ) );
  AND2X1_RVT U807 ( .A1(n75), .A2(n52), .Y(\ab[0][16] ) );
  AND2X1_RVT U808 ( .A1(n75), .A2(n49), .Y(\ab[0][15] ) );
  AND2X1_RVT U809 ( .A1(n75), .A2(n46), .Y(\ab[0][14] ) );
  AND2X1_RVT U810 ( .A1(n75), .A2(n43), .Y(\ab[0][13] ) );
  AND2X1_RVT U811 ( .A1(n75), .A2(n40), .Y(\ab[0][12] ) );
  AND2X1_RVT U812 ( .A1(n75), .A2(n37), .Y(\ab[0][11] ) );
  AND2X1_RVT U813 ( .A1(n75), .A2(n34), .Y(\ab[0][10] ) );
  AND2X1_RVT U814 ( .A1(n75), .A2(n4), .Y(PRODUCT[0]) );
endmodule


module fpu_DW_div_uns_2 ( a, b, quotient, remainder, divide_by_0 );
  input [46:0] a;
  input [23:0] b;
  output [46:0] quotient;
  output [23:0] remainder;
  output divide_by_0;
  wire   \u_div/SumTmp[1][1] , \u_div/SumTmp[1][2] , \u_div/SumTmp[1][3] ,
         \u_div/SumTmp[1][4] , \u_div/SumTmp[1][5] , \u_div/SumTmp[1][6] ,
         \u_div/SumTmp[1][7] , \u_div/SumTmp[1][8] , \u_div/SumTmp[1][9] ,
         \u_div/SumTmp[1][10] , \u_div/SumTmp[1][11] , \u_div/SumTmp[1][12] ,
         \u_div/SumTmp[1][13] , \u_div/SumTmp[1][14] , \u_div/SumTmp[1][15] ,
         \u_div/SumTmp[1][16] , \u_div/SumTmp[1][17] , \u_div/SumTmp[1][18] ,
         \u_div/SumTmp[1][19] , \u_div/SumTmp[1][20] , \u_div/SumTmp[1][21] ,
         \u_div/SumTmp[1][22] , \u_div/SumTmp[1][23] , \u_div/SumTmp[2][1] ,
         \u_div/SumTmp[2][2] , \u_div/SumTmp[2][3] , \u_div/SumTmp[2][4] ,
         \u_div/SumTmp[2][5] , \u_div/SumTmp[2][6] , \u_div/SumTmp[2][7] ,
         \u_div/SumTmp[2][8] , \u_div/SumTmp[2][9] , \u_div/SumTmp[2][10] ,
         \u_div/SumTmp[2][11] , \u_div/SumTmp[2][12] , \u_div/SumTmp[2][13] ,
         \u_div/SumTmp[2][14] , \u_div/SumTmp[2][15] , \u_div/SumTmp[2][16] ,
         \u_div/SumTmp[2][17] , \u_div/SumTmp[2][18] , \u_div/SumTmp[2][19] ,
         \u_div/SumTmp[2][20] , \u_div/SumTmp[2][21] , \u_div/SumTmp[2][22] ,
         \u_div/SumTmp[2][23] , \u_div/SumTmp[3][1] , \u_div/SumTmp[3][2] ,
         \u_div/SumTmp[3][3] , \u_div/SumTmp[3][4] , \u_div/SumTmp[3][5] ,
         \u_div/SumTmp[3][6] , \u_div/SumTmp[3][7] , \u_div/SumTmp[3][8] ,
         \u_div/SumTmp[3][9] , \u_div/SumTmp[3][10] , \u_div/SumTmp[3][11] ,
         \u_div/SumTmp[3][12] , \u_div/SumTmp[3][13] , \u_div/SumTmp[3][14] ,
         \u_div/SumTmp[3][15] , \u_div/SumTmp[3][16] , \u_div/SumTmp[3][17] ,
         \u_div/SumTmp[3][18] , \u_div/SumTmp[3][19] , \u_div/SumTmp[3][20] ,
         \u_div/SumTmp[3][21] , \u_div/SumTmp[3][22] , \u_div/SumTmp[3][23] ,
         \u_div/SumTmp[4][1] , \u_div/SumTmp[4][2] , \u_div/SumTmp[4][3] ,
         \u_div/SumTmp[4][4] , \u_div/SumTmp[4][5] , \u_div/SumTmp[4][6] ,
         \u_div/SumTmp[4][7] , \u_div/SumTmp[4][8] , \u_div/SumTmp[4][9] ,
         \u_div/SumTmp[4][10] , \u_div/SumTmp[4][11] , \u_div/SumTmp[4][12] ,
         \u_div/SumTmp[4][13] , \u_div/SumTmp[4][14] , \u_div/SumTmp[4][15] ,
         \u_div/SumTmp[4][16] , \u_div/SumTmp[4][17] , \u_div/SumTmp[4][18] ,
         \u_div/SumTmp[4][19] , \u_div/SumTmp[4][20] , \u_div/SumTmp[4][21] ,
         \u_div/SumTmp[5][0] , \u_div/SumTmp[5][1] , \u_div/SumTmp[5][2] ,
         \u_div/SumTmp[5][3] , \u_div/SumTmp[5][5] , \u_div/SumTmp[5][6] ,
         \u_div/SumTmp[5][7] , \u_div/SumTmp[5][8] , \u_div/SumTmp[5][9] ,
         \u_div/SumTmp[5][23] , \u_div/SumTmp[6][0] , \u_div/SumTmp[6][1] ,
         \u_div/SumTmp[6][2] , \u_div/SumTmp[6][3] , \u_div/SumTmp[6][4] ,
         \u_div/SumTmp[6][5] , \u_div/SumTmp[6][6] , \u_div/SumTmp[6][10] ,
         \u_div/SumTmp[6][11] , \u_div/SumTmp[6][12] , \u_div/SumTmp[6][13] ,
         \u_div/SumTmp[6][14] , \u_div/SumTmp[6][15] , \u_div/SumTmp[6][16] ,
         \u_div/SumTmp[6][17] , \u_div/SumTmp[6][18] , \u_div/SumTmp[6][19] ,
         \u_div/SumTmp[6][20] , \u_div/SumTmp[6][21] , \u_div/SumTmp[6][22] ,
         \u_div/SumTmp[6][23] , \u_div/SumTmp[7][0] , \u_div/SumTmp[7][1] ,
         \u_div/SumTmp[7][2] , \u_div/SumTmp[7][3] , \u_div/SumTmp[7][4] ,
         \u_div/SumTmp[7][5] , \u_div/SumTmp[7][6] , \u_div/SumTmp[7][7] ,
         \u_div/SumTmp[7][9] , \u_div/SumTmp[7][10] , \u_div/SumTmp[7][11] ,
         \u_div/SumTmp[7][12] , \u_div/SumTmp[7][13] , \u_div/SumTmp[7][14] ,
         \u_div/SumTmp[7][15] , \u_div/SumTmp[7][16] , \u_div/SumTmp[7][17] ,
         \u_div/SumTmp[7][19] , \u_div/SumTmp[8][0] , \u_div/SumTmp[8][1] ,
         \u_div/SumTmp[8][2] , \u_div/SumTmp[8][3] , \u_div/SumTmp[8][4] ,
         \u_div/SumTmp[8][5] , \u_div/SumTmp[8][7] , \u_div/SumTmp[8][8] ,
         \u_div/SumTmp[8][9] , \u_div/SumTmp[8][10] , \u_div/SumTmp[8][11] ,
         \u_div/SumTmp[8][12] , \u_div/SumTmp[8][13] , \u_div/SumTmp[8][14] ,
         \u_div/SumTmp[8][15] , \u_div/SumTmp[8][16] , \u_div/SumTmp[8][17] ,
         \u_div/SumTmp[8][18] , \u_div/SumTmp[8][20] , \u_div/SumTmp[8][21] ,
         \u_div/SumTmp[8][22] , \u_div/SumTmp[9][0] , \u_div/SumTmp[9][1] ,
         \u_div/SumTmp[9][2] , \u_div/SumTmp[9][3] , \u_div/SumTmp[9][4] ,
         \u_div/SumTmp[9][19] , \u_div/SumTmp[9][20] , \u_div/SumTmp[9][21] ,
         \u_div/SumTmp[9][22] , \u_div/SumTmp[9][23] , \u_div/SumTmp[10][1] ,
         \u_div/SumTmp[10][2] , \u_div/SumTmp[10][3] , \u_div/SumTmp[10][5] ,
         \u_div/SumTmp[10][6] , \u_div/SumTmp[10][7] , \u_div/SumTmp[10][8] ,
         \u_div/SumTmp[10][9] , \u_div/SumTmp[10][10] , \u_div/SumTmp[10][11] ,
         \u_div/SumTmp[11][0] , \u_div/SumTmp[11][1] , \u_div/SumTmp[11][2] ,
         \u_div/SumTmp[11][3] , \u_div/SumTmp[11][4] , \u_div/SumTmp[11][5] ,
         \u_div/SumTmp[11][6] , \u_div/SumTmp[11][7] , \u_div/SumTmp[11][8] ,
         \u_div/SumTmp[11][9] , \u_div/SumTmp[11][10] , \u_div/SumTmp[11][12] ,
         \u_div/SumTmp[11][13] , \u_div/SumTmp[11][14] ,
         \u_div/SumTmp[11][15] , \u_div/SumTmp[11][16] ,
         \u_div/SumTmp[11][17] , \u_div/SumTmp[11][18] ,
         \u_div/SumTmp[11][19] , \u_div/SumTmp[11][20] ,
         \u_div/SumTmp[11][21] , \u_div/SumTmp[12][0] , \u_div/SumTmp[12][1] ,
         \u_div/SumTmp[12][2] , \u_div/SumTmp[12][3] , \u_div/SumTmp[12][4] ,
         \u_div/SumTmp[12][5] , \u_div/SumTmp[12][6] , \u_div/SumTmp[12][7] ,
         \u_div/SumTmp[12][8] , \u_div/SumTmp[12][9] , \u_div/SumTmp[12][10] ,
         \u_div/SumTmp[12][11] , \u_div/SumTmp[12][12] ,
         \u_div/SumTmp[12][13] , \u_div/SumTmp[12][14] ,
         \u_div/SumTmp[12][15] , \u_div/SumTmp[12][17] ,
         \u_div/SumTmp[12][18] , \u_div/SumTmp[12][19] ,
         \u_div/SumTmp[12][20] , \u_div/SumTmp[12][22] , \u_div/SumTmp[13][0] ,
         \u_div/SumTmp[13][1] , \u_div/SumTmp[13][2] , \u_div/SumTmp[13][3] ,
         \u_div/SumTmp[13][4] , \u_div/SumTmp[13][5] , \u_div/SumTmp[13][6] ,
         \u_div/SumTmp[13][7] , \u_div/SumTmp[13][8] , \u_div/SumTmp[13][9] ,
         \u_div/SumTmp[13][10] , \u_div/SumTmp[13][11] ,
         \u_div/SumTmp[13][13] , \u_div/SumTmp[13][14] ,
         \u_div/SumTmp[13][15] , \u_div/SumTmp[13][16] ,
         \u_div/SumTmp[13][17] , \u_div/SumTmp[13][18] ,
         \u_div/SumTmp[13][19] , \u_div/SumTmp[13][21] ,
         \u_div/SumTmp[13][22] , \u_div/SumTmp[13][23] , \u_div/SumTmp[14][0] ,
         \u_div/SumTmp[14][1] , \u_div/SumTmp[14][2] , \u_div/SumTmp[14][3] ,
         \u_div/SumTmp[14][4] , \u_div/SumTmp[14][5] , \u_div/SumTmp[14][6] ,
         \u_div/SumTmp[14][7] , \u_div/SumTmp[14][8] , \u_div/SumTmp[14][9] ,
         \u_div/SumTmp[14][10] , \u_div/SumTmp[14][11] ,
         \u_div/SumTmp[14][20] , \u_div/SumTmp[14][21] ,
         \u_div/SumTmp[14][22] , \u_div/SumTmp[14][23] , \u_div/SumTmp[15][0] ,
         \u_div/SumTmp[15][1] , \u_div/SumTmp[15][2] , \u_div/SumTmp[15][3] ,
         \u_div/SumTmp[15][4] , \u_div/SumTmp[15][5] , \u_div/SumTmp[15][6] ,
         \u_div/SumTmp[15][7] , \u_div/SumTmp[15][8] , \u_div/SumTmp[15][9] ,
         \u_div/SumTmp[15][10] , \u_div/SumTmp[15][12] ,
         \u_div/SumTmp[15][13] , \u_div/SumTmp[16][0] , \u_div/SumTmp[16][14] ,
         \u_div/SumTmp[16][15] , \u_div/SumTmp[16][17] ,
         \u_div/SumTmp[16][18] , \u_div/SumTmp[16][19] ,
         \u_div/SumTmp[16][20] , \u_div/SumTmp[16][21] ,
         \u_div/SumTmp[16][22] , \u_div/SumTmp[17][1] , \u_div/SumTmp[17][2] ,
         \u_div/SumTmp[17][3] , \u_div/SumTmp[17][4] , \u_div/SumTmp[17][5] ,
         \u_div/SumTmp[17][6] , \u_div/SumTmp[17][7] , \u_div/SumTmp[17][8] ,
         \u_div/SumTmp[17][9] , \u_div/SumTmp[17][10] , \u_div/SumTmp[17][11] ,
         \u_div/SumTmp[17][12] , \u_div/SumTmp[17][13] ,
         \u_div/SumTmp[17][14] , \u_div/SumTmp[17][15] ,
         \u_div/SumTmp[17][16] , \u_div/SumTmp[17][17] ,
         \u_div/SumTmp[17][18] , \u_div/SumTmp[17][19] , \u_div/SumTmp[18][0] ,
         \u_div/SumTmp[18][1] , \u_div/SumTmp[18][2] , \u_div/SumTmp[18][3] ,
         \u_div/SumTmp[18][4] , \u_div/SumTmp[18][5] , \u_div/SumTmp[18][6] ,
         \u_div/SumTmp[18][7] , \u_div/SumTmp[18][8] , \u_div/SumTmp[18][9] ,
         \u_div/SumTmp[18][10] , \u_div/SumTmp[18][11] ,
         \u_div/SumTmp[18][12] , \u_div/SumTmp[18][13] ,
         \u_div/SumTmp[18][14] , \u_div/SumTmp[18][15] ,
         \u_div/SumTmp[18][16] , \u_div/SumTmp[19][0] , \u_div/SumTmp[19][1] ,
         \u_div/SumTmp[19][2] , \u_div/SumTmp[19][3] , \u_div/SumTmp[19][4] ,
         \u_div/SumTmp[19][5] , \u_div/SumTmp[19][6] , \u_div/SumTmp[19][7] ,
         \u_div/SumTmp[19][8] , \u_div/SumTmp[19][9] , \u_div/SumTmp[19][10] ,
         \u_div/SumTmp[19][11] , \u_div/SumTmp[19][12] ,
         \u_div/SumTmp[19][13] , \u_div/SumTmp[19][14] ,
         \u_div/SumTmp[19][15] , \u_div/SumTmp[20][0] , \u_div/SumTmp[20][1] ,
         \u_div/SumTmp[20][2] , \u_div/SumTmp[20][3] , \u_div/SumTmp[20][4] ,
         \u_div/SumTmp[20][5] , \u_div/SumTmp[20][6] , \u_div/SumTmp[20][7] ,
         \u_div/SumTmp[20][8] , \u_div/SumTmp[20][9] , \u_div/SumTmp[20][10] ,
         \u_div/SumTmp[20][11] , \u_div/SumTmp[20][17] ,
         \u_div/SumTmp[20][18] , \u_div/SumTmp[20][19] ,
         \u_div/SumTmp[20][20] , \u_div/SumTmp[20][21] ,
         \u_div/SumTmp[20][22] , \u_div/SumTmp[21][0] , \u_div/SumTmp[21][1] ,
         \u_div/SumTmp[21][2] , \u_div/SumTmp[21][3] , \u_div/SumTmp[21][4] ,
         \u_div/SumTmp[21][5] , \u_div/SumTmp[21][12] , \u_div/SumTmp[21][13] ,
         \u_div/SumTmp[21][14] , \u_div/SumTmp[21][15] ,
         \u_div/SumTmp[21][16] , \u_div/SumTmp[21][17] ,
         \u_div/SumTmp[21][18] , \u_div/SumTmp[21][19] ,
         \u_div/SumTmp[21][20] , \u_div/SumTmp[21][21] ,
         \u_div/SumTmp[21][22] , \u_div/SumTmp[21][23] , \u_div/SumTmp[22][0] ,
         \u_div/SumTmp[22][1] , \u_div/SumTmp[22][2] , \u_div/SumTmp[22][3] ,
         \u_div/SumTmp[22][6] , \u_div/SumTmp[22][7] , \u_div/SumTmp[22][8] ,
         \u_div/SumTmp[22][9] , \u_div/SumTmp[22][10] , \u_div/SumTmp[22][11] ,
         \u_div/SumTmp[22][12] , \u_div/SumTmp[22][13] ,
         \u_div/SumTmp[22][14] , \u_div/SumTmp[22][15] ,
         \u_div/SumTmp[22][16] , \u_div/SumTmp[22][17] ,
         \u_div/SumTmp[22][18] , \u_div/SumTmp[22][19] ,
         \u_div/SumTmp[22][20] , \u_div/SumTmp[22][21] ,
         \u_div/SumTmp[22][22] , \u_div/SumTmp[22][23] , \u_div/SumTmp[23][1] ,
         \u_div/SumTmp[23][2] , \u_div/SumTmp[23][3] , \u_div/SumTmp[23][4] ,
         \u_div/SumTmp[23][5] , \u_div/SumTmp[23][6] , \u_div/SumTmp[23][7] ,
         \u_div/SumTmp[23][8] , \u_div/SumTmp[23][9] , \u_div/SumTmp[23][10] ,
         \u_div/SumTmp[23][11] , \u_div/SumTmp[23][12] ,
         \u_div/SumTmp[23][13] , \u_div/SumTmp[23][14] ,
         \u_div/SumTmp[23][15] , \u_div/SumTmp[23][16] ,
         \u_div/SumTmp[23][17] , \u_div/SumTmp[23][18] ,
         \u_div/SumTmp[23][19] , \u_div/SumTmp[23][20] ,
         \u_div/SumTmp[23][21] , \u_div/SumTmp[24][1] , \u_div/SumTmp[24][2] ,
         \u_div/SumTmp[24][3] , \u_div/SumTmp[24][4] , \u_div/SumTmp[24][5] ,
         \u_div/SumTmp[24][6] , \u_div/SumTmp[24][7] , \u_div/SumTmp[24][8] ,
         \u_div/SumTmp[24][9] , \u_div/SumTmp[24][10] , \u_div/SumTmp[24][11] ,
         \u_div/SumTmp[24][12] , \u_div/SumTmp[24][13] ,
         \u_div/SumTmp[24][22] , \u_div/SumTmp[25][1] , \u_div/SumTmp[25][2] ,
         \u_div/SumTmp[25][3] , \u_div/SumTmp[25][4] , \u_div/SumTmp[25][5] ,
         \u_div/SumTmp[25][6] , \u_div/SumTmp[25][7] , \u_div/SumTmp[25][8] ,
         \u_div/SumTmp[26][1] , \u_div/SumTmp[26][2] , \u_div/SumTmp[26][3] ,
         \u_div/SumTmp[26][4] , \u_div/SumTmp[26][5] , \u_div/SumTmp[26][6] ,
         \u_div/SumTmp[26][7] , \u_div/SumTmp[26][9] , \u_div/SumTmp[26][10] ,
         \u_div/SumTmp[27][1] , \u_div/SumTmp[27][2] , \u_div/SumTmp[27][3] ,
         \u_div/SumTmp[27][4] , \u_div/SumTmp[27][5] , \u_div/SumTmp[27][6] ,
         \u_div/SumTmp[27][7] , \u_div/SumTmp[27][8] , \u_div/SumTmp[27][9] ,
         \u_div/SumTmp[27][11] , \u_div/SumTmp[27][12] ,
         \u_div/SumTmp[27][13] , \u_div/SumTmp[27][14] ,
         \u_div/SumTmp[27][15] , \u_div/SumTmp[27][16] ,
         \u_div/SumTmp[27][17] , \u_div/SumTmp[27][18] ,
         \u_div/SumTmp[27][19] , \u_div/SumTmp[28][10] ,
         \u_div/SumTmp[28][11] , \u_div/SumTmp[28][12] ,
         \u_div/SumTmp[28][13] , \u_div/SumTmp[28][14] ,
         \u_div/SumTmp[28][15] , \u_div/SumTmp[28][16] ,
         \u_div/SumTmp[28][17] , \u_div/SumTmp[28][18] , \u_div/SumTmp[29][1] ,
         \u_div/SumTmp[29][2] , \u_div/SumTmp[29][3] , \u_div/SumTmp[29][4] ,
         \u_div/SumTmp[29][5] , \u_div/SumTmp[29][6] , \u_div/SumTmp[29][7] ,
         \u_div/SumTmp[29][8] , \u_div/SumTmp[29][9] , \u_div/SumTmp[29][10] ,
         \u_div/SumTmp[29][11] , \u_div/SumTmp[29][12] ,
         \u_div/SumTmp[29][13] , \u_div/SumTmp[29][14] ,
         \u_div/SumTmp[29][15] , \u_div/SumTmp[29][16] , \u_div/SumTmp[30][1] ,
         \u_div/SumTmp[30][2] , \u_div/SumTmp[30][3] , \u_div/SumTmp[30][4] ,
         \u_div/SumTmp[30][5] , \u_div/SumTmp[30][6] , \u_div/SumTmp[30][7] ,
         \u_div/SumTmp[30][8] , \u_div/SumTmp[30][9] , \u_div/SumTmp[30][10] ,
         \u_div/SumTmp[30][11] , \u_div/SumTmp[30][12] ,
         \u_div/SumTmp[30][13] , \u_div/SumTmp[30][14] , \u_div/SumTmp[31][1] ,
         \u_div/SumTmp[31][2] , \u_div/SumTmp[31][3] , \u_div/SumTmp[31][4] ,
         \u_div/SumTmp[31][5] , \u_div/SumTmp[31][6] , \u_div/SumTmp[31][7] ,
         \u_div/SumTmp[31][8] , \u_div/SumTmp[31][9] , \u_div/SumTmp[31][10] ,
         \u_div/SumTmp[31][11] , \u_div/SumTmp[31][12] ,
         \u_div/SumTmp[31][13] , \u_div/SumTmp[31][15] , \u_div/SumTmp[32][1] ,
         \u_div/SumTmp[32][2] , \u_div/SumTmp[32][3] , \u_div/SumTmp[32][4] ,
         \u_div/SumTmp[32][5] , \u_div/SumTmp[32][6] , \u_div/SumTmp[32][7] ,
         \u_div/SumTmp[32][8] , \u_div/SumTmp[32][9] , \u_div/SumTmp[32][10] ,
         \u_div/SumTmp[33][1] , \u_div/SumTmp[33][2] , \u_div/SumTmp[33][3] ,
         \u_div/SumTmp[33][4] , \u_div/SumTmp[33][5] , \u_div/SumTmp[33][6] ,
         \u_div/SumTmp[33][7] , \u_div/SumTmp[33][8] , \u_div/SumTmp[33][9] ,
         \u_div/SumTmp[33][11] , \u_div/SumTmp[33][12] ,
         \u_div/SumTmp[33][13] , \u_div/SumTmp[34][1] , \u_div/SumTmp[34][2] ,
         \u_div/SumTmp[34][3] , \u_div/SumTmp[34][4] , \u_div/SumTmp[34][10] ,
         \u_div/SumTmp[34][11] , \u_div/SumTmp[34][12] , \u_div/SumTmp[35][1] ,
         \u_div/SumTmp[35][2] , \u_div/SumTmp[35][3] , \u_div/SumTmp[35][5] ,
         \u_div/SumTmp[35][6] , \u_div/SumTmp[35][7] , \u_div/SumTmp[35][8] ,
         \u_div/SumTmp[35][9] , \u_div/SumTmp[35][10] , \u_div/SumTmp[35][11] ,
         \u_div/SumTmp[36][1] , \u_div/SumTmp[36][2] , \u_div/SumTmp[36][4] ,
         \u_div/SumTmp[36][5] , \u_div/SumTmp[36][6] , \u_div/SumTmp[36][7] ,
         \u_div/SumTmp[36][8] , \u_div/SumTmp[36][9] , \u_div/SumTmp[36][10] ,
         \u_div/SumTmp[37][3] , \u_div/SumTmp[37][4] , \u_div/SumTmp[37][5] ,
         \u_div/SumTmp[37][6] , \u_div/SumTmp[37][7] , \u_div/SumTmp[37][8] ,
         \u_div/SumTmp[37][9] , \u_div/SumTmp[38][2] , \u_div/SumTmp[38][3] ,
         \u_div/SumTmp[38][4] , \u_div/SumTmp[38][5] , \u_div/SumTmp[38][6] ,
         \u_div/SumTmp[39][1] , \u_div/SumTmp[39][2] , \u_div/SumTmp[39][3] ,
         \u_div/SumTmp[39][4] , \u_div/SumTmp[39][5] , \u_div/SumTmp[40][1] ,
         \u_div/SumTmp[40][2] , \u_div/SumTmp[40][3] , \u_div/SumTmp[40][4] ,
         \u_div/SumTmp[40][5] , \u_div/SumTmp[41][1] , \u_div/SumTmp[41][2] ,
         \u_div/SumTmp[41][3] , \u_div/SumTmp[41][4] , \u_div/SumTmp[42][1] ,
         \u_div/SumTmp[42][2] , \u_div/SumTmp[42][3] , \u_div/SumTmp[44][1] ,
         \u_div/SumTmp[44][2] , \u_div/SumTmp[45][1] , \u_div/CryTmp[0][2] ,
         \u_div/CryTmp[0][3] , \u_div/CryTmp[0][4] , \u_div/CryTmp[0][5] ,
         \u_div/CryTmp[0][6] , \u_div/CryTmp[0][7] , \u_div/CryTmp[0][8] ,
         \u_div/CryTmp[0][9] , \u_div/CryTmp[0][10] , \u_div/CryTmp[0][11] ,
         \u_div/CryTmp[0][12] , \u_div/CryTmp[0][13] , \u_div/CryTmp[0][14] ,
         \u_div/CryTmp[0][15] , \u_div/CryTmp[0][16] , \u_div/CryTmp[0][17] ,
         \u_div/CryTmp[0][18] , \u_div/CryTmp[0][19] , \u_div/CryTmp[0][20] ,
         \u_div/CryTmp[0][21] , \u_div/CryTmp[0][22] , \u_div/CryTmp[0][23] ,
         \u_div/CryTmp[0][24] , \u_div/CryTmp[1][2] , \u_div/CryTmp[1][3] ,
         \u_div/CryTmp[1][4] , \u_div/CryTmp[1][5] , \u_div/CryTmp[1][6] ,
         \u_div/CryTmp[1][7] , \u_div/CryTmp[1][8] , \u_div/CryTmp[1][9] ,
         \u_div/CryTmp[1][10] , \u_div/CryTmp[1][11] , \u_div/CryTmp[1][12] ,
         \u_div/CryTmp[1][13] , \u_div/CryTmp[1][14] , \u_div/CryTmp[1][15] ,
         \u_div/CryTmp[1][16] , \u_div/CryTmp[1][17] , \u_div/CryTmp[1][18] ,
         \u_div/CryTmp[1][19] , \u_div/CryTmp[1][20] , \u_div/CryTmp[1][21] ,
         \u_div/CryTmp[1][22] , \u_div/CryTmp[1][23] , \u_div/CryTmp[1][24] ,
         \u_div/CryTmp[2][2] , \u_div/CryTmp[2][3] , \u_div/CryTmp[2][4] ,
         \u_div/CryTmp[2][5] , \u_div/CryTmp[2][6] , \u_div/CryTmp[2][7] ,
         \u_div/CryTmp[2][8] , \u_div/CryTmp[2][9] , \u_div/CryTmp[2][10] ,
         \u_div/CryTmp[2][11] , \u_div/CryTmp[2][12] , \u_div/CryTmp[2][13] ,
         \u_div/CryTmp[2][14] , \u_div/CryTmp[2][15] , \u_div/CryTmp[2][16] ,
         \u_div/CryTmp[2][17] , \u_div/CryTmp[2][18] , \u_div/CryTmp[2][19] ,
         \u_div/CryTmp[2][20] , \u_div/CryTmp[2][21] , \u_div/CryTmp[2][22] ,
         \u_div/CryTmp[2][23] , \u_div/CryTmp[2][24] , \u_div/CryTmp[5][23] ,
         \u_div/CryTmp[5][24] , \u_div/CryTmp[6][11] , \u_div/CryTmp[6][12] ,
         \u_div/CryTmp[6][13] , \u_div/CryTmp[6][14] , \u_div/CryTmp[6][15] ,
         \u_div/CryTmp[6][16] , \u_div/CryTmp[6][17] , \u_div/CryTmp[6][18] ,
         \u_div/CryTmp[6][19] , \u_div/CryTmp[6][20] , \u_div/CryTmp[6][21] ,
         \u_div/CryTmp[6][22] , \u_div/CryTmp[6][23] , \u_div/CryTmp[6][24] ,
         \u_div/CryTmp[7][9] , \u_div/CryTmp[7][10] , \u_div/CryTmp[7][11] ,
         \u_div/CryTmp[7][12] , \u_div/CryTmp[7][13] , \u_div/CryTmp[7][14] ,
         \u_div/CryTmp[7][15] , \u_div/CryTmp[7][16] , \u_div/CryTmp[7][17] ,
         \u_div/CryTmp[7][18] , \u_div/CryTmp[8][24] , \u_div/CryTmp[9][20] ,
         \u_div/CryTmp[9][21] , \u_div/CryTmp[9][22] , \u_div/CryTmp[9][23] ,
         \u_div/CryTmp[9][24] , \u_div/CryTmp[11][1] , \u_div/CryTmp[12][24] ,
         \u_div/CryTmp[13][21] , \u_div/CryTmp[13][22] ,
         \u_div/CryTmp[13][23] , \u_div/CryTmp[13][24] ,
         \u_div/CryTmp[14][21] , \u_div/CryTmp[14][22] ,
         \u_div/CryTmp[14][23] , \u_div/CryTmp[14][24] ,
         \u_div/CryTmp[16][24] , \u_div/CryTmp[20][24] ,
         \u_div/CryTmp[21][13] , \u_div/CryTmp[21][14] ,
         \u_div/CryTmp[21][15] , \u_div/CryTmp[21][16] ,
         \u_div/CryTmp[21][17] , \u_div/CryTmp[21][18] ,
         \u_div/CryTmp[21][19] , \u_div/CryTmp[21][20] ,
         \u_div/CryTmp[21][21] , \u_div/CryTmp[21][22] ,
         \u_div/CryTmp[21][23] , \u_div/CryTmp[21][24] , \u_div/CryTmp[22][1] ,
         \u_div/CryTmp[22][6] , \u_div/CryTmp[22][7] , \u_div/CryTmp[22][8] ,
         \u_div/CryTmp[22][9] , \u_div/CryTmp[22][10] , \u_div/CryTmp[22][11] ,
         \u_div/CryTmp[22][12] , \u_div/CryTmp[22][13] ,
         \u_div/CryTmp[22][14] , \u_div/CryTmp[22][15] ,
         \u_div/CryTmp[22][16] , \u_div/CryTmp[24][23] ,
         \u_div/CryTmp[27][11] , \u_div/CryTmp[27][12] ,
         \u_div/CryTmp[27][13] , \u_div/CryTmp[27][14] ,
         \u_div/CryTmp[27][15] , \u_div/CryTmp[27][16] ,
         \u_div/CryTmp[27][17] , \u_div/CryTmp[27][18] ,
         \u_div/CryTmp[27][19] , \u_div/CryTmp[27][20] ,
         \u_div/CryTmp[28][11] , \u_div/CryTmp[28][12] ,
         \u_div/CryTmp[28][13] , \u_div/CryTmp[28][14] ,
         \u_div/CryTmp[28][15] , \u_div/CryTmp[28][16] ,
         \u_div/CryTmp[28][17] , \u_div/CryTmp[28][18] ,
         \u_div/CryTmp[28][19] , \u_div/CryTmp[31][15] ,
         \u_div/CryTmp[31][16] , \u_div/CryTmp[33][11] ,
         \u_div/CryTmp[33][12] , \u_div/CryTmp[33][13] ,
         \u_div/CryTmp[33][14] , \u_div/CryTmp[34][11] ,
         \u_div/CryTmp[34][12] , \u_div/CryTmp[34][13] , \u_div/CryTmp[35][5] ,
         \u_div/CryTmp[35][6] , \u_div/CryTmp[35][7] , \u_div/CryTmp[35][8] ,
         \u_div/CryTmp[35][9] , \u_div/CryTmp[35][10] , \u_div/CryTmp[35][11] ,
         \u_div/CryTmp[35][12] , \u_div/CryTmp[36][4] , \u_div/CryTmp[36][5] ,
         \u_div/CryTmp[36][6] , \u_div/CryTmp[36][7] , \u_div/CryTmp[36][8] ,
         \u_div/CryTmp[36][9] , \u_div/CryTmp[36][10] , \u_div/CryTmp[36][11] ,
         \u_div/CryTmp[37][4] , \u_div/CryTmp[37][5] , \u_div/CryTmp[37][6] ,
         \u_div/CryTmp[37][7] , \u_div/CryTmp[37][8] , \u_div/CryTmp[37][9] ,
         \u_div/CryTmp[37][10] , \u_div/CryTmp[40][7] , \u_div/CryTmp[41][6] ,
         \u_div/CryTmp[42][5] , \u_div/CryTmp[45][1] , \u_div/CryTmp[45][2] ,
         \u_div/PartRem[1][1] , \u_div/PartRem[1][2] , \u_div/PartRem[1][3] ,
         \u_div/PartRem[1][4] , \u_div/PartRem[1][5] , \u_div/PartRem[1][6] ,
         \u_div/PartRem[1][7] , \u_div/PartRem[1][8] , \u_div/PartRem[1][9] ,
         \u_div/PartRem[1][10] , \u_div/PartRem[1][11] ,
         \u_div/PartRem[1][12] , \u_div/PartRem[1][13] ,
         \u_div/PartRem[1][14] , \u_div/PartRem[1][15] ,
         \u_div/PartRem[1][16] , \u_div/PartRem[1][17] ,
         \u_div/PartRem[1][18] , \u_div/PartRem[1][19] ,
         \u_div/PartRem[1][20] , \u_div/PartRem[1][21] ,
         \u_div/PartRem[1][22] , \u_div/PartRem[1][23] ,
         \u_div/PartRem[1][24] , \u_div/PartRem[2][1] , \u_div/PartRem[2][2] ,
         \u_div/PartRem[2][3] , \u_div/PartRem[2][4] , \u_div/PartRem[2][5] ,
         \u_div/PartRem[2][6] , \u_div/PartRem[2][7] , \u_div/PartRem[2][9] ,
         \u_div/PartRem[2][10] , \u_div/PartRem[2][13] ,
         \u_div/PartRem[2][14] , \u_div/PartRem[2][15] ,
         \u_div/PartRem[2][16] , \u_div/PartRem[2][17] ,
         \u_div/PartRem[2][18] , \u_div/PartRem[2][19] ,
         \u_div/PartRem[2][20] , \u_div/PartRem[2][21] ,
         \u_div/PartRem[2][22] , \u_div/PartRem[2][23] ,
         \u_div/PartRem[2][24] , \u_div/PartRem[3][1] , \u_div/PartRem[3][2] ,
         \u_div/PartRem[3][3] , \u_div/PartRem[3][4] , \u_div/PartRem[3][5] ,
         \u_div/PartRem[3][6] , \u_div/PartRem[3][7] , \u_div/PartRem[3][8] ,
         \u_div/PartRem[3][9] , \u_div/PartRem[3][10] , \u_div/PartRem[3][12] ,
         \u_div/PartRem[3][13] , \u_div/PartRem[3][14] ,
         \u_div/PartRem[3][15] , \u_div/PartRem[3][16] ,
         \u_div/PartRem[3][17] , \u_div/PartRem[3][18] ,
         \u_div/PartRem[3][19] , \u_div/PartRem[3][20] ,
         \u_div/PartRem[3][21] , \u_div/PartRem[3][22] ,
         \u_div/PartRem[3][23] , \u_div/PartRem[3][24] ,
         \u_div/PartRem[5][24] , \u_div/PartRem[6][6] , \u_div/PartRem[6][24] ,
         \u_div/PartRem[7][6] , \u_div/PartRem[7][10] , \u_div/PartRem[7][11] ,
         \u_div/PartRem[7][12] , \u_div/PartRem[7][13] ,
         \u_div/PartRem[7][14] , \u_div/PartRem[7][15] ,
         \u_div/PartRem[7][16] , \u_div/PartRem[7][17] ,
         \u_div/PartRem[7][18] , \u_div/PartRem[7][19] ,
         \u_div/PartRem[7][20] , \u_div/PartRem[7][21] ,
         \u_div/PartRem[7][22] , \u_div/PartRem[7][23] ,
         \u_div/PartRem[7][24] , \u_div/PartRem[8][9] , \u_div/PartRem[8][10] ,
         \u_div/PartRem[8][12] , \u_div/PartRem[8][13] ,
         \u_div/PartRem[8][14] , \u_div/PartRem[8][15] ,
         \u_div/PartRem[8][16] , \u_div/PartRem[8][17] ,
         \u_div/PartRem[8][18] , \u_div/PartRem[9][10] ,
         \u_div/PartRem[9][24] , \u_div/PartRem[10][19] ,
         \u_div/PartRem[10][20] , \u_div/PartRem[10][21] ,
         \u_div/PartRem[10][22] , \u_div/PartRem[10][23] ,
         \u_div/PartRem[10][24] , \u_div/PartRem[13][24] ,
         \u_div/PartRem[14][21] , \u_div/PartRem[14][22] ,
         \u_div/PartRem[14][23] , \u_div/PartRem[14][24] ,
         \u_div/PartRem[15][20] , \u_div/PartRem[15][21] ,
         \u_div/PartRem[15][22] , \u_div/PartRem[15][23] ,
         \u_div/PartRem[15][24] , \u_div/PartRem[17][24] ,
         \u_div/PartRem[21][24] , \u_div/PartRem[22][12] ,
         \u_div/PartRem[22][13] , \u_div/PartRem[22][14] ,
         \u_div/PartRem[22][15] , \u_div/PartRem[22][16] ,
         \u_div/PartRem[22][17] , \u_div/PartRem[22][18] ,
         \u_div/PartRem[22][19] , \u_div/PartRem[22][20] ,
         \u_div/PartRem[22][21] , \u_div/PartRem[22][22] ,
         \u_div/PartRem[22][23] , \u_div/PartRem[22][24] ,
         \u_div/PartRem[23][6] , \u_div/PartRem[23][7] ,
         \u_div/PartRem[23][8] , \u_div/PartRem[23][9] ,
         \u_div/PartRem[23][10] , \u_div/PartRem[23][11] ,
         \u_div/PartRem[23][12] , \u_div/PartRem[23][13] ,
         \u_div/PartRem[23][14] , \u_div/PartRem[23][15] ,
         \u_div/PartRem[23][16] , \u_div/PartRem[23][23] ,
         \u_div/PartRem[25][22] , \u_div/PartRem[28][11] ,
         \u_div/PartRem[28][12] , \u_div/PartRem[28][13] ,
         \u_div/PartRem[28][14] , \u_div/PartRem[28][15] ,
         \u_div/PartRem[28][16] , \u_div/PartRem[28][17] ,
         \u_div/PartRem[28][18] , \u_div/PartRem[28][19] ,
         \u_div/PartRem[29][10] , \u_div/PartRem[29][11] ,
         \u_div/PartRem[29][12] , \u_div/PartRem[29][13] ,
         \u_div/PartRem[29][14] , \u_div/PartRem[29][15] ,
         \u_div/PartRem[29][16] , \u_div/PartRem[29][17] ,
         \u_div/PartRem[29][18] , \u_div/PartRem[32][15] ,
         \u_div/PartRem[34][11] , \u_div/PartRem[34][12] ,
         \u_div/PartRem[34][13] , \u_div/PartRem[35][8] ,
         \u_div/PartRem[35][10] , \u_div/PartRem[35][11] ,
         \u_div/PartRem[35][12] , \u_div/PartRem[36][3] ,
         \u_div/PartRem[36][5] , \u_div/PartRem[36][6] ,
         \u_div/PartRem[36][7] , \u_div/PartRem[36][8] ,
         \u_div/PartRem[36][9] , \u_div/PartRem[36][10] ,
         \u_div/PartRem[36][11] , \u_div/PartRem[37][4] ,
         \u_div/PartRem[37][5] , \u_div/PartRem[37][6] ,
         \u_div/PartRem[37][7] , \u_div/PartRem[37][8] ,
         \u_div/PartRem[37][9] , \u_div/PartRem[37][10] ,
         \u_div/PartRem[38][4] , \u_div/PartRem[38][5] ,
         \u_div/PartRem[38][6] , \u_div/PartRem[38][7] ,
         \u_div/PartRem[38][8] , \u_div/PartRem[38][9] ,
         \u_div/PartRem[39][2] , \u_div/PartRem[39][5] ,
         \u_div/PartRem[39][6] , \u_div/PartRem[46][1] , net31320, net31310,
         net31303, net31297, net31295, net31294, net31292, net31291, net31287,
         net31281, net31276, net31273, net31272, net31271, net31270, net31261,
         net31255, net31250, net31244, net31243, net31242, net31213, net31212,
         net31211, net31209, net31208, net31207, net31206, net31205, net31204,
         net31203, net31202, net31201, net31200, net31198, net31197, net31196,
         net31195, net31194, net31193, net31192, net31191, net31190, net31189,
         net31188, net31186, net31185, net31184, net31183, net31182, net31181,
         net31180, net31179, net31178, net31177, net31176, net31175, net31173,
         net31172, net31171, net31170, net31168, net31165, net31164, net31163,
         net31162, net31161, net31160, net31158, net31157, net31156, net31155,
         net31154, net31153, net31150, net31149, net31148, net31147, net31146,
         net31145, net31144, net31142, net31141, net31140, net31139, net31138,
         net31137, net31134, net31133, net31132, net31131, net31130, net31129,
         net31128, net31127, net31125, net31124, net31123, net31122, net31121,
         net31120, net31117, net31116, net31115, net31113, net31112, net31111,
         net31110, net31109, net31105, net31104, net31103, net31099, net31098,
         net31097, net31096, net31093, net31092, net31091, net31090, net31088,
         net31086, net31085, net31084, net31080, net31079, net31078, net31077,
         net31076, net31075, net31073, net31072, net31071, net31070, net31068,
         net31066, net31065, net31064, net31063, net31058, net31057, net31056,
         net31055, net31054, net31053, net31051, net31050, net31049, net31048,
         net31044, net31043, net31042, net31041, net31038, net31036, net31035,
         net31034, net31033, net31032, net31031, net31029, net31028, net31027,
         net31026, net31025, net31024, net31022, net31021, net31020, net31019,
         net31016, net31015, net31013, net31012, net31011, net31010, net31009,
         net31008, net31006, net31005, net31004, net31003, net31002, net31001,
         net30999, net30998, net30997, net30996, net30993, net30992, net30991,
         net30989, net30988, net30987, net30986, net30985, net30984, net30981,
         net30980, net30979, net30978, net30977, net30975, net30974, net30973,
         net30972, net30968, net30967, net30966, net30965, net30963, net30962,
         net30961, net30960, net30959, net30957, net30955, net30954, net30953,
         net30952, net30951, net30946, net30945, net30944, net30943, net30942,
         net30941, net30940, net30939, net30938, net30937, net30936, net30935,
         net30934, net30933, net30931, net30930, net30929, net30928, net30927,
         net30926, net30925, net30924, net30923, net30922, net30921, net30920,
         net30919, net30916, net30915, net30914, net30913, net30912, net30911,
         net30910, net30909, net30907, net30906, net30905, net30904, net30903,
         net30902, net30899, net30893, net30892, net30890, net30889, net30888,
         net30885, net30884, net30883, net30882, net30881, net30879, net30876,
         net30875, net30873, net30871, net30870, net30869, net30868, net30867,
         net30866, net30865, net30864, net30863, net30853, net30838, net30837,
         net30836, net30835, net30834, net30833, net30831, net30830, net30828,
         net30827, net30825, net30821, net30820, net30819, net30816, net30807,
         net30801, net30794, net30791, net30790, net30789, net30788, net30787,
         net30786, net30785, net30783, net30782, net30780, net30779, net30777,
         net30773, net30772, net30771, net30758, net30748, net30744, net30743,
         net30742, net30741, net30740, net30739, net30738, net30737, net30733,
         net30732, net30731, net30729, net30728, net30724, net30723, net30702,
         net30696, net30695, net30694, net30693, net30692, net30691, net30690,
         net30689, net30687, net30686, net30683, net30681, net30680, net30677,
         net30676, net30675, net30666, net30664, net30663, net30661, net30660,
         net30659, net30658, net30657, net30656, net30655, net30654, net30653,
         net30645, net30644, net30643, net30642, net30641, net30639, net30638,
         net30636, net30635, net30634, net30633, net30632, net30629, net30628,
         net30627, net30626, net30625, net30624, net30623, net30622, net30621,
         net30620, net30613, net30606, net30603, net30599, net30598, net30597,
         net30596, net30595, net30594, net30593, net30591, net30590, net30588,
         net30587, net30586, net30585, net30584, net30583, net30572, net30571,
         net30570, net30569, net30568, net30567, net30566, net30565, net30564,
         net30563, net30562, net30560, net30559, net30556, net30555, net30554,
         net30551, net30549, net30548, net30547, net30546, net30545, net30543,
         net30542, net30540, net30539, net30538, net30537, net30536, net30535,
         net30534, net30533, net30532, net30531, net30530, net30529, net30528,
         net30527, net30526, net30512, net30509, net30508, net30507, net30506,
         net30501, net30500, net30499, net30498, net30497, net30495, net30494,
         net30492, net30491, net30490, net30489, net30488, net30487, net30478,
         net30476, net30475, net30474, net30473, net30472, net30471, net30468,
         net30466, net30465, net30464, net30462, net30461, net30458, net30456,
         net30455, net30453, net30452, net30451, net30448, net30446, net30445,
         net30443, net30442, net30441, net30435, net30433, net30432, net30431,
         net30426, net30422, net30421, net30416, net30414, net30412, net30411,
         net30406, net30404, net30402, net30401, net30398, net30397, net30394,
         net30392, net30391, net30386, net30384, net30382, net30381, net30376,
         net30374, net30372, net30371, net30366, net30364, net30362, net30361,
         net30358, net30357, net30356, net30354, net30352, net30351, net30346,
         net30344, net30342, net30341, net30336, net30335, net30334, net30332,
         net30331, net30322, net30318, net30317, net30314, net30313, net30312,
         net30311, net30308, net30307, net30306, net30305, net30304, net30301,
         net30300, net30299, net30298, net30297, net30296, net30293, net30291,
         net30290, net30289, net30288, net30287, net30286, net30271, net30270,
         net30267, net30266, net30265, net30264, net30260, net30256, net30255,
         net30254, net30252, net30251, net30249, net30248, net30247, net30245,
         net30223, net30219, net30218, net30217, net30216, net30211, net30210,
         net30208, net30207, net30206, net30204, net30203, net30202, net30200,
         net30199, net30187, net30186, net30185, net30184, net30183, net30182,
         net30181, net30180, net30178, net30177, net30161, net30159, net30158,
         net30157, net30150, net30146, net30144, net30143, net30142, net30135,
         net30130, net30124, net30123, net30122, net30121, net30119, net30118,
         net30117, net30099, net30098, net30087, net30086, net30085, net30081,
         net30080, net30079, net30074, net30072, net30071, net30070, net30069,
         net30068, net30067, net30066, net30065, net30064, net30063, net30053,
         net30051, net30050, net30049, net30048, net30047, net30036, net30033,
         net30022, net30015, net30013, net30012, net29982, net29981, net29980,
         net29979, net29978, net29977, net29976, net29975, net29974, net29956,
         net29944, net29942, net29940, net29939, net29937, net29936, net29935,
         net29934, net29933, net29932, net29931, net29921, net29899, net29885,
         net29874, net29873, net29872, net29862, net29854, net29852, net29846,
         net29844, net29843, net29841, net29837, net29822, net29821, net29820,
         net29819, net29818, net29817, net29816, net29815, net29801, net29796,
         net29795, net29782, net29779, net29778, net29755, net29753, net29752,
         net29751, net29750, net29749, net29748, net29747, net29746, net29744,
         net29743, net29742, net29741, net29737, net29733, net29732, net29731,
         net29730, net29729, net29728, net29727, net29726, net29711, net29710,
         net29709, net29708, net29702, net29698, net29685, net29684, net29683,
         net29682, net29681, net29680, net29676, net29674, net29672, net29671,
         net29670, net29669, net29668, net29667, net29666, net29665, net29664,
         net29663, net29662, net29661, net29658, net29656, net29655, net29654,
         net29653, net29649, net29648, net29647, net29646, net29637, net29636,
         net29635, net29632, net29631, net29628, net29624, net29623, net29622,
         net29619, net29618, net29617, net29616, net29615, net29614, net29613,
         net29612, net29606, net29599, net29598, net31434, net31466, net31482,
         net31498, net31514, net31530, net31562, net31578, net31594, net31610,
         net31626, net31642, net31658, net31674, net31706, net31722, net31738,
         net31770, net31786, net31802, net31800, net31822, net31814, net31828,
         net31826, net31846, net31844, net31856, net31854, net31874, net31872,
         net31884, net31882, net31902, net31896, net31914, net31912, net31910,
         net31930, net31922, net31940, net31938, net31952, net31950, net31964,
         net31962, net31960, net31974, net31972, net31986, net31984, net31982,
         net32002, net31998, net32016, net32014, net32012, net32032, net32024,
         net32046, net32044, net32042, net32068, net32066, net32078, net32076,
         net32092, net32090, net32088, net32106, net32104, net32118, net32116,
         net32130, net32128, net32144, net32142, net32140, net32156, net32154,
         net32168, net32166, net32186, net32178, net32200, net32198, net32196,
         net32212, net32210, net32226, net32224, net32222, net32242, net32234,
         net32254, net32252, net32250, net32272, net32264, net32284, net32282,
         net32280, net32302, net32300, net32314, net32312, net32310, net32326,
         net32324, net32338, net32336, net32334, net32354, net32352, net32368,
         net32366, net32364, net32362, net32386, net32384, net32382, net32408,
         net32406, net32506, net32520, net32518, net32530, net32538, net32536,
         net32544, net32542, net32550, net32548, net32554, net32560, net32568,
         net32566, net32580, net32578, net32592, net32590, net32598, net32596,
         net32610, net32608, net32616, net32624, net32620,
         \*cell*33666/net34045 , \*cell*33669/net34055 ,
         \*cell*33672/net34065 , \*cell*33675/net34075 ,
         \*cell*33681/net34095 , \*cell*33684/net34105 ,
         \*cell*33687/net34115 , \*cell*33690/net34125 ,
         \*cell*33693/net34135 , \*cell*33696/net34145 ,
         \*cell*33702/net34165 , \*cell*33717/net34215 ,
         \*cell*33720/net34225 , \*cell*33723/net34235 ,
         \*cell*33726/net34245 , net37169, net37184, net37220, net37219,
         net37224, net37228, net37229, net37231, net37242, net37244, net37246,
         net37247, net37248, net37249, net37251, net37252, net37253, net37254,
         net37256, net37261, net37263, net37556, net37563, net37567, net37570,
         net37577, net37581, net37584, net37585, net37854, net38272, net38274,
         net38337, net38341, net38342, net38343, net38350, net39870, net39869,
         net39874, net39872, net40084, net40598, net40656, net40724, net40721,
         net40720, net40719, net40718, net40717, net40783, net41046, net41045,
         net41415, net41435, net42034, net42041, net42040, net42357, net42365,
         net42408, net42398, net42397, net42523, net42520, net42519, net42517,
         net42516, net42515, net42514, net42512, net42548, net42939, net42938,
         net43355, net43354, net43819, net43885, net43884, net44064, net44063,
         net44395, net44394, net44464, net44466, net44755, net44969, net44967,
         net45002, net45007, net45183, net45229, net45228, net45257, net45288,
         net45295, net45541, net45604, net45603, net45602, net45601, net45600,
         net45599, net45597, net45594, net45592, net45588, net45587, net45585,
         net45584, net45583, net45582, net45581, net45654, net45678, net45677,
         net45671, net45669, net45665, net45737, net46142, net46238, net46242,
         net46241, net46343, net46421, net46550, net46608, net46688, net46768,
         net46859, net46962, net46961, net47679, net47688, net47690, net47709,
         net47716, net47718, net47729, net47816, net47979, net47978, net48342,
         net48341, net48340, net48339, net48385, net48384, net48534, net48533,
         net48639, net48638, net48659, net48658, net48671, net48670, net48759,
         net48758, net49055, net49113, net49112, net49213, net49212, net49211,
         net49255, net49254, net49281, net49280, net49311, net49310, net49309,
         net49601, net49608, net49612, net49611, net49616, net49626, net49625,
         net49675, net49674, net49679, net49678, net50050, net50049, net50177,
         net50176, net50182, net50186, net50185, net50339, net50471, net50470,
         net50727, net50726, net50743, net50742, net51612, net51611, net51994,
         net52000, net52003, net52013, net52012, net52520, net52534, net52536,
         net52890, net52992, net52991, \u_div/SumTmp[8][6] ,
         \u_div/SumTmp[8][23] , \u_div/SumTmp[7][8] , \u_div/SumTmp[7][23] ,
         \u_div/SumTmp[7][22] , \u_div/SumTmp[7][21] , \u_div/SumTmp[7][20] ,
         \u_div/SumTmp[6][9] , \u_div/SumTmp[6][8] , \u_div/SumTmp[6][7] ,
         \u_div/SumTmp[5][4] , \u_div/SumTmp[5][22] , \u_div/SumTmp[5][21] ,
         \u_div/SumTmp[5][20] , \u_div/SumTmp[5][19] , \u_div/SumTmp[5][18] ,
         \u_div/SumTmp[5][17] , \u_div/SumTmp[5][16] , \u_div/SumTmp[5][15] ,
         \u_div/SumTmp[5][14] , \u_div/SumTmp[5][13] , \u_div/SumTmp[5][12] ,
         \u_div/SumTmp[5][11] , \u_div/SumTmp[5][10] , \u_div/SumTmp[4][23] ,
         \u_div/SumTmp[4][22] , \u_div/PartRem[9][6] , \u_div/PartRem[9][23] ,
         \u_div/PartRem[9][22] , \u_div/PartRem[9][21] ,
         \u_div/PartRem[9][20] , \u_div/PartRem[8][8] , \u_div/PartRem[8][6] ,
         \u_div/PartRem[8][5] , \u_div/PartRem[8][4] , \u_div/PartRem[8][3] ,
         \u_div/PartRem[8][2] , \u_div/PartRem[8][24] , \u_div/PartRem[8][23] ,
         \u_div/PartRem[8][22] , \u_div/PartRem[8][1] , \u_div/PartRem[8][19] ,
         \u_div/PartRem[7][9] , \u_div/PartRem[7][8] , \u_div/PartRem[7][7] ,
         \u_div/PartRem[7][5] , \u_div/PartRem[7][4] , \u_div/PartRem[7][3] ,
         \u_div/PartRem[7][2] , \u_div/PartRem[7][1] , \u_div/PartRem[6][5] ,
         \u_div/PartRem[6][4] , \u_div/PartRem[6][3] , \u_div/PartRem[6][2] ,
         \u_div/PartRem[6][21] , \u_div/PartRem[6][20] , \u_div/PartRem[6][1] ,
         \u_div/PartRem[6][19] , \u_div/PartRem[6][18] ,
         \u_div/PartRem[6][17] , \u_div/PartRem[6][16] ,
         \u_div/PartRem[6][15] , \u_div/PartRem[6][14] ,
         \u_div/PartRem[6][13] , \u_div/PartRem[6][12] ,
         \u_div/PartRem[6][11] , \u_div/PartRem[5][9] , \u_div/PartRem[5][8] ,
         \u_div/PartRem[5][6] , \u_div/PartRem[5][5] , \u_div/PartRem[5][4] ,
         \u_div/PartRem[5][3] , \u_div/PartRem[5][2] , \u_div/PartRem[5][21] ,
         \u_div/PartRem[5][20] , \u_div/PartRem[5][1] , \u_div/PartRem[5][19] ,
         \u_div/PartRem[5][18] , \u_div/PartRem[5][17] ,
         \u_div/PartRem[5][16] , \u_div/PartRem[5][15] ,
         \u_div/PartRem[5][14] , \u_div/PartRem[5][13] ,
         \u_div/PartRem[5][12] , \u_div/PartRem[5][11] ,
         \u_div/PartRem[5][10] , \u_div/PartRem[4][9] , \u_div/PartRem[4][8] ,
         \u_div/PartRem[4][7] , \u_div/PartRem[4][6] , \u_div/PartRem[4][5] ,
         \u_div/PartRem[4][4] , \u_div/PartRem[4][3] , \u_div/PartRem[4][2] ,
         \u_div/PartRem[4][24] , \u_div/PartRem[4][22] ,
         \u_div/PartRem[4][21] , \u_div/PartRem[4][20] , \u_div/PartRem[4][1] ,
         \u_div/PartRem[4][19] , \u_div/PartRem[4][18] ,
         \u_div/PartRem[4][17] , \u_div/PartRem[4][16] ,
         \u_div/PartRem[4][15] , \u_div/PartRem[4][14] ,
         \u_div/PartRem[4][13] , \u_div/PartRem[4][12] ,
         \u_div/PartRem[4][11] , \u_div/PartRem[4][10] , \u_div/CryTmp[8][23] ,
         \u_div/CryTmp[8][22] , \u_div/CryTmp[8][21] , \u_div/CryTmp[8][20] ,
         \u_div/CryTmp[7][8] , \u_div/CryTmp[7][7] , \u_div/CryTmp[7][6] ,
         \u_div/CryTmp[7][5] , \u_div/CryTmp[7][4] , \u_div/CryTmp[7][3] ,
         \u_div/CryTmp[7][2] , \u_div/CryTmp[7][24] , \u_div/CryTmp[7][23] ,
         \u_div/CryTmp[7][22] , \u_div/CryTmp[7][21] , \u_div/CryTmp[7][20] ,
         \u_div/CryTmp[7][19] , \u_div/CryTmp[6][9] , \u_div/CryTmp[6][8] ,
         \u_div/CryTmp[6][7] , \u_div/CryTmp[6][6] , \u_div/CryTmp[6][5] ,
         \u_div/CryTmp[6][4] , \u_div/CryTmp[6][3] , \u_div/CryTmp[6][2] ,
         \u_div/CryTmp[6][10] , \u_div/CryTmp[5][9] , \u_div/CryTmp[5][8] ,
         \u_div/CryTmp[5][7] , \u_div/CryTmp[5][6] , \u_div/CryTmp[5][5] ,
         \u_div/CryTmp[5][4] , \u_div/CryTmp[5][3] , \u_div/CryTmp[5][2] ,
         \u_div/CryTmp[5][22] , \u_div/CryTmp[5][21] , \u_div/CryTmp[5][20] ,
         \u_div/CryTmp[5][19] , \u_div/CryTmp[5][18] , \u_div/CryTmp[5][17] ,
         \u_div/CryTmp[5][16] , \u_div/CryTmp[5][15] , \u_div/CryTmp[5][14] ,
         \u_div/CryTmp[5][13] , \u_div/CryTmp[5][12] , \u_div/CryTmp[5][11] ,
         \u_div/CryTmp[5][10] , \u_div/CryTmp[4][9] , \u_div/CryTmp[4][8] ,
         \u_div/CryTmp[4][7] , \u_div/CryTmp[4][6] , \u_div/CryTmp[4][5] ,
         \u_div/CryTmp[4][4] , \u_div/CryTmp[4][3] , \u_div/CryTmp[4][2] ,
         \u_div/CryTmp[4][24] , \u_div/CryTmp[4][23] , \u_div/CryTmp[4][22] ,
         \u_div/CryTmp[4][21] , \u_div/CryTmp[4][20] , \u_div/CryTmp[4][19] ,
         \u_div/CryTmp[4][18] , \u_div/CryTmp[4][17] , \u_div/CryTmp[4][16] ,
         \u_div/CryTmp[4][15] , \u_div/CryTmp[4][14] , \u_div/CryTmp[4][13] ,
         \u_div/CryTmp[4][12] , \u_div/CryTmp[4][11] , \u_div/CryTmp[4][10] ,
         \u_div/CryTmp[3][9] , \u_div/CryTmp[3][8] , \u_div/CryTmp[3][7] ,
         \u_div/CryTmp[3][6] , \u_div/CryTmp[3][5] , \u_div/CryTmp[3][4] ,
         \u_div/CryTmp[3][3] , \u_div/CryTmp[3][2] , \u_div/CryTmp[3][24] ,
         \u_div/CryTmp[3][23] , \u_div/CryTmp[3][22] , \u_div/CryTmp[3][21] ,
         \u_div/CryTmp[3][20] , \u_div/CryTmp[3][19] , \u_div/CryTmp[3][18] ,
         \u_div/CryTmp[3][17] , \u_div/CryTmp[3][16] , \u_div/CryTmp[3][15] ,
         \u_div/CryTmp[3][14] , \u_div/CryTmp[3][13] , \u_div/CryTmp[3][12] ,
         \u_div/CryTmp[3][11] , \u_div/CryTmp[3][10] , net38347, net29611,
         net29609, net29605, net29604, net29603, net29602, net29600,
         \u_div/SumTmp[9][9] , \u_div/SumTmp[9][8] , \u_div/SumTmp[9][7] ,
         \u_div/SumTmp[9][6] , \u_div/SumTmp[9][5] , \u_div/SumTmp[9][18] ,
         \u_div/SumTmp[9][17] , \u_div/SumTmp[9][16] , \u_div/SumTmp[9][15] ,
         \u_div/SumTmp[9][14] , \u_div/SumTmp[9][13] , \u_div/SumTmp[9][12] ,
         \u_div/SumTmp[9][11] , \u_div/SumTmp[9][10] , \u_div/SumTmp[8][19] ,
         \u_div/SumTmp[10][4] , \u_div/SumTmp[10][23] , \u_div/SumTmp[10][22] ,
         \u_div/SumTmp[10][21] , \u_div/SumTmp[10][20] ,
         \u_div/SumTmp[10][19] , \u_div/SumTmp[10][18] ,
         \u_div/SumTmp[10][17] , \u_div/SumTmp[10][16] , \u_div/PartRem[9][9] ,
         \u_div/PartRem[9][8] , \u_div/PartRem[9][7] , \u_div/PartRem[9][5] ,
         \u_div/PartRem[9][4] , \u_div/PartRem[9][3] , \u_div/PartRem[9][2] ,
         \u_div/PartRem[9][1] , \u_div/PartRem[9][19] , \u_div/PartRem[9][18] ,
         \u_div/PartRem[9][17] , \u_div/PartRem[9][16] ,
         \u_div/PartRem[9][15] , \u_div/PartRem[9][14] ,
         \u_div/PartRem[9][13] , \u_div/PartRem[9][12] ,
         \u_div/PartRem[9][11] , \u_div/PartRem[8][20] ,
         \u_div/PartRem[11][24] , \u_div/PartRem[11][23] ,
         \u_div/PartRem[11][22] , \u_div/PartRem[11][21] ,
         \u_div/PartRem[11][20] , \u_div/PartRem[11][19] ,
         \u_div/PartRem[11][18] , \u_div/PartRem[11][17] ,
         \u_div/PartRem[11][16] , \u_div/PartRem[10][9] ,
         \u_div/PartRem[10][8] , \u_div/PartRem[10][7] ,
         \u_div/PartRem[10][6] , \u_div/PartRem[10][5] ,
         \u_div/PartRem[10][4] , \u_div/PartRem[10][3] ,
         \u_div/PartRem[10][2] , \u_div/PartRem[10][1] ,
         \u_div/PartRem[10][18] , \u_div/PartRem[10][17] ,
         \u_div/PartRem[10][16] , \u_div/PartRem[10][15] ,
         \u_div/PartRem[10][14] , \u_div/PartRem[10][13] ,
         \u_div/PartRem[10][12] , \u_div/PartRem[10][11] ,
         \u_div/PartRem[10][10] , \u_div/CryTmp[9][9] , \u_div/CryTmp[9][8] ,
         \u_div/CryTmp[9][7] , \u_div/CryTmp[9][6] , \u_div/CryTmp[9][5] ,
         \u_div/CryTmp[9][4] , \u_div/CryTmp[9][3] , \u_div/CryTmp[9][2] ,
         \u_div/CryTmp[9][19] , \u_div/CryTmp[9][18] , \u_div/CryTmp[9][17] ,
         \u_div/CryTmp[9][16] , \u_div/CryTmp[9][15] , \u_div/CryTmp[9][14] ,
         \u_div/CryTmp[9][13] , \u_div/CryTmp[9][12] , \u_div/CryTmp[9][11] ,
         \u_div/CryTmp[9][10] , \u_div/CryTmp[8][9] , \u_div/CryTmp[8][8] ,
         \u_div/CryTmp[8][7] , \u_div/CryTmp[8][6] , \u_div/CryTmp[8][5] ,
         \u_div/CryTmp[8][4] , \u_div/CryTmp[8][3] , \u_div/CryTmp[8][2] ,
         \u_div/CryTmp[8][19] , \u_div/CryTmp[8][18] , \u_div/CryTmp[8][17] ,
         \u_div/CryTmp[8][16] , \u_div/CryTmp[8][15] , \u_div/CryTmp[8][14] ,
         \u_div/CryTmp[8][13] , \u_div/CryTmp[8][12] , \u_div/CryTmp[8][11] ,
         \u_div/CryTmp[8][10] , \u_div/CryTmp[10][24] , \u_div/CryTmp[10][23] ,
         \u_div/CryTmp[10][22] , \u_div/CryTmp[10][21] ,
         \u_div/CryTmp[10][20] , \u_div/CryTmp[10][19] ,
         \u_div/CryTmp[10][18] , \u_div/CryTmp[10][17] , net31102, net30932,
         net30901, net30900, net30898, net30897, net30896, net30895, net30891,
         net30862, net30861, net30860, net30859, net30858, net30857, net30856,
         net30855, net30849, net30848, net30846, net30845, net30843, net30842,
         net30477, net30467, net30457, net30447, net30428, net30427, net30418,
         net30417, net30408, net30407, net30388, net30387, net30378, net30377,
         net30368, net30367, net30348, net30347, net30338, net30337, net29946,
         net29945, net29798, net29797, net29740, net29739, net29738, net29633,
         net29601, \u_div/SumTmp[14][19] , \u_div/SumTmp[14][18] ,
         \u_div/SumTmp[14][17] , \u_div/SumTmp[14][16] ,
         \u_div/SumTmp[14][15] , \u_div/SumTmp[14][14] ,
         \u_div/SumTmp[14][13] , \u_div/SumTmp[14][12] ,
         \u_div/SumTmp[13][20] , \u_div/SumTmp[13][12] ,
         \u_div/SumTmp[12][23] , \u_div/SumTmp[12][21] ,
         \u_div/SumTmp[12][16] , \u_div/SumTmp[11][23] ,
         \u_div/SumTmp[11][22] , \u_div/SumTmp[11][11] ,
         \u_div/SumTmp[10][15] , \u_div/SumTmp[10][14] ,
         \u_div/SumTmp[10][13] , \u_div/SumTmp[10][12] ,
         \u_div/PartRem[15][9] , \u_div/PartRem[15][8] ,
         \u_div/PartRem[15][7] , \u_div/PartRem[15][6] ,
         \u_div/PartRem[15][5] , \u_div/PartRem[15][4] ,
         \u_div/PartRem[15][3] , \u_div/PartRem[15][2] ,
         \u_div/PartRem[15][1] , \u_div/PartRem[15][19] ,
         \u_div/PartRem[15][18] , \u_div/PartRem[15][17] ,
         \u_div/PartRem[15][16] , \u_div/PartRem[15][15] ,
         \u_div/PartRem[15][14] , \u_div/PartRem[15][13] ,
         \u_div/PartRem[15][11] , \u_div/PartRem[15][10] ,
         \u_div/PartRem[14][9] , \u_div/PartRem[14][8] ,
         \u_div/PartRem[14][7] , \u_div/PartRem[14][6] ,
         \u_div/PartRem[14][5] , \u_div/PartRem[14][4] ,
         \u_div/PartRem[14][3] , \u_div/PartRem[14][2] ,
         \u_div/PartRem[14][20] , \u_div/PartRem[14][1] ,
         \u_div/PartRem[14][19] , \u_div/PartRem[14][18] ,
         \u_div/PartRem[14][17] , \u_div/PartRem[14][16] ,
         \u_div/PartRem[14][15] , \u_div/PartRem[14][14] ,
         \u_div/PartRem[14][13] , \u_div/PartRem[14][12] ,
         \u_div/PartRem[14][11] , \u_div/PartRem[14][10] ,
         \u_div/PartRem[13][9] , \u_div/PartRem[13][8] ,
         \u_div/PartRem[13][7] , \u_div/PartRem[13][6] ,
         \u_div/PartRem[13][5] , \u_div/PartRem[13][4] ,
         \u_div/PartRem[13][3] , \u_div/PartRem[13][2] ,
         \u_div/PartRem[13][23] , \u_div/PartRem[13][22] ,
         \u_div/PartRem[13][21] , \u_div/PartRem[13][20] ,
         \u_div/PartRem[13][1] , \u_div/PartRem[13][19] ,
         \u_div/PartRem[13][18] , \u_div/PartRem[13][17] ,
         \u_div/PartRem[13][16] , \u_div/PartRem[13][15] ,
         \u_div/PartRem[13][14] , \u_div/PartRem[13][13] ,
         \u_div/PartRem[13][12] , \u_div/PartRem[13][11] ,
         \u_div/PartRem[13][10] , \u_div/PartRem[12][9] ,
         \u_div/PartRem[12][8] , \u_div/PartRem[12][7] ,
         \u_div/PartRem[12][6] , \u_div/PartRem[12][5] ,
         \u_div/PartRem[12][4] , \u_div/PartRem[12][3] ,
         \u_div/PartRem[12][2] , \u_div/PartRem[12][24] ,
         \u_div/PartRem[12][23] , \u_div/PartRem[12][22] ,
         \u_div/PartRem[12][21] , \u_div/PartRem[12][20] ,
         \u_div/PartRem[12][1] , \u_div/PartRem[12][19] ,
         \u_div/PartRem[12][18] , \u_div/PartRem[12][17] ,
         \u_div/PartRem[12][16] , \u_div/PartRem[12][15] ,
         \u_div/PartRem[12][14] , \u_div/PartRem[12][13] ,
         \u_div/PartRem[12][12] , \u_div/PartRem[12][10] ,
         \u_div/PartRem[11][9] , \u_div/PartRem[11][8] ,
         \u_div/PartRem[11][7] , \u_div/PartRem[11][6] ,
         \u_div/PartRem[11][5] , \u_div/PartRem[11][4] ,
         \u_div/PartRem[11][3] , \u_div/PartRem[11][2] ,
         \u_div/PartRem[11][1] , \u_div/PartRem[11][15] ,
         \u_div/PartRem[11][14] , \u_div/PartRem[11][13] ,
         \u_div/PartRem[11][11] , \u_div/PartRem[11][10] ,
         \u_div/CryTmp[14][9] , \u_div/CryTmp[14][8] , \u_div/CryTmp[14][7] ,
         \u_div/CryTmp[14][6] , \u_div/CryTmp[14][5] , \u_div/CryTmp[14][4] ,
         \u_div/CryTmp[14][3] , \u_div/CryTmp[14][2] , \u_div/CryTmp[14][20] ,
         \u_div/CryTmp[14][19] , \u_div/CryTmp[14][18] ,
         \u_div/CryTmp[14][17] , \u_div/CryTmp[14][16] ,
         \u_div/CryTmp[14][15] , \u_div/CryTmp[14][14] ,
         \u_div/CryTmp[14][13] , \u_div/CryTmp[14][12] ,
         \u_div/CryTmp[14][11] , \u_div/CryTmp[14][10] , \u_div/CryTmp[13][9] ,
         \u_div/CryTmp[13][8] , \u_div/CryTmp[13][7] , \u_div/CryTmp[13][6] ,
         \u_div/CryTmp[13][5] , \u_div/CryTmp[13][4] , \u_div/CryTmp[13][3] ,
         \u_div/CryTmp[13][2] , \u_div/CryTmp[13][20] , \u_div/CryTmp[13][19] ,
         \u_div/CryTmp[13][18] , \u_div/CryTmp[13][17] ,
         \u_div/CryTmp[13][16] , \u_div/CryTmp[13][15] ,
         \u_div/CryTmp[13][14] , \u_div/CryTmp[13][13] ,
         \u_div/CryTmp[13][12] , \u_div/CryTmp[13][11] ,
         \u_div/CryTmp[13][10] , \u_div/CryTmp[12][9] , \u_div/CryTmp[12][8] ,
         \u_div/CryTmp[12][7] , \u_div/CryTmp[12][6] , \u_div/CryTmp[12][5] ,
         \u_div/CryTmp[12][4] , \u_div/CryTmp[12][3] , \u_div/CryTmp[12][2] ,
         \u_div/CryTmp[12][23] , \u_div/CryTmp[12][22] ,
         \u_div/CryTmp[12][21] , \u_div/CryTmp[12][20] ,
         \u_div/CryTmp[12][19] , \u_div/CryTmp[12][18] ,
         \u_div/CryTmp[12][17] , \u_div/CryTmp[12][16] ,
         \u_div/CryTmp[12][15] , \u_div/CryTmp[12][14] ,
         \u_div/CryTmp[12][13] , \u_div/CryTmp[12][12] ,
         \u_div/CryTmp[12][11] , \u_div/CryTmp[12][10] , \u_div/CryTmp[11][9] ,
         \u_div/CryTmp[11][8] , \u_div/CryTmp[11][7] , \u_div/CryTmp[11][6] ,
         \u_div/CryTmp[11][5] , \u_div/CryTmp[11][4] , \u_div/CryTmp[11][3] ,
         \u_div/CryTmp[11][2] , \u_div/CryTmp[11][24] , \u_div/CryTmp[11][23] ,
         \u_div/CryTmp[11][22] , \u_div/CryTmp[11][21] ,
         \u_div/CryTmp[11][20] , \u_div/CryTmp[11][19] ,
         \u_div/CryTmp[11][18] , \u_div/CryTmp[11][17] ,
         \u_div/CryTmp[11][16] , \u_div/CryTmp[11][15] ,
         \u_div/CryTmp[11][14] , \u_div/CryTmp[11][13] ,
         \u_div/CryTmp[11][12] , \u_div/CryTmp[11][11] ,
         \u_div/CryTmp[11][10] , \u_div/CryTmp[10][9] , \u_div/CryTmp[10][8] ,
         \u_div/CryTmp[10][7] , \u_div/CryTmp[10][6] , \u_div/CryTmp[10][5] ,
         \u_div/CryTmp[10][4] , \u_div/CryTmp[10][3] , \u_div/CryTmp[10][2] ,
         \u_div/CryTmp[10][16] , \u_div/CryTmp[10][15] ,
         \u_div/CryTmp[10][14] , \u_div/CryTmp[10][13] ,
         \u_div/CryTmp[10][12] , \u_div/CryTmp[10][11] ,
         \u_div/CryTmp[10][10] , net49094, net46895, net46752, net45940,
         net45939, net42406, net42405, net38336, net31106, net30948, net30947,
         net30841, net30806, net30805, net30803, net30802, net30800, net30799,
         net30798, net30797, net30796, net30795, net30768, net30767, net30766,
         net30765, net30764, net30763, net30762, net30761, net30757, net30755,
         net30708, \u_div/SumTmp[16][9] , \u_div/SumTmp[16][8] ,
         \u_div/SumTmp[16][7] , \u_div/SumTmp[16][6] , \u_div/SumTmp[16][5] ,
         \u_div/SumTmp[16][4] , \u_div/SumTmp[16][3] , \u_div/SumTmp[16][2] ,
         \u_div/SumTmp[16][23] , \u_div/SumTmp[16][1] , \u_div/SumTmp[16][16] ,
         \u_div/SumTmp[16][13] , \u_div/SumTmp[16][12] ,
         \u_div/SumTmp[16][11] , \u_div/SumTmp[16][10] ,
         \u_div/SumTmp[15][23] , \u_div/SumTmp[15][22] ,
         \u_div/SumTmp[15][21] , \u_div/SumTmp[15][20] ,
         \u_div/SumTmp[15][19] , \u_div/SumTmp[15][18] ,
         \u_div/SumTmp[15][17] , \u_div/SumTmp[15][16] ,
         \u_div/SumTmp[15][15] , \u_div/SumTmp[15][14] ,
         \u_div/SumTmp[15][11] , \u_div/PartRem[17][9] ,
         \u_div/PartRem[17][8] , \u_div/PartRem[17][7] ,
         \u_div/PartRem[17][6] , \u_div/PartRem[17][5] ,
         \u_div/PartRem[17][4] , \u_div/PartRem[17][3] ,
         \u_div/PartRem[17][2] , \u_div/PartRem[17][23] ,
         \u_div/PartRem[17][22] , \u_div/PartRem[17][21] ,
         \u_div/PartRem[17][20] , \u_div/PartRem[17][19] ,
         \u_div/PartRem[17][18] , \u_div/PartRem[17][17] ,
         \u_div/PartRem[17][16] , \u_div/PartRem[17][15] ,
         \u_div/PartRem[17][14] , \u_div/PartRem[17][13] ,
         \u_div/PartRem[17][12] , \u_div/PartRem[17][11] ,
         \u_div/PartRem[17][10] , \u_div/PartRem[16][9] ,
         \u_div/PartRem[16][8] , \u_div/PartRem[16][7] ,
         \u_div/PartRem[16][6] , \u_div/PartRem[16][5] ,
         \u_div/PartRem[16][4] , \u_div/PartRem[16][3] ,
         \u_div/PartRem[16][2] , \u_div/PartRem[16][24] ,
         \u_div/PartRem[16][23] , \u_div/PartRem[16][22] ,
         \u_div/PartRem[16][21] , \u_div/PartRem[16][20] ,
         \u_div/PartRem[16][1] , \u_div/PartRem[16][19] ,
         \u_div/PartRem[16][18] , \u_div/PartRem[16][17] ,
         \u_div/PartRem[16][16] , \u_div/PartRem[16][15] ,
         \u_div/PartRem[16][14] , \u_div/PartRem[16][13] ,
         \u_div/PartRem[16][12] , \u_div/PartRem[16][11] ,
         \u_div/PartRem[16][10] , \u_div/PartRem[15][12] ,
         \u_div/CryTmp[16][9] , \u_div/CryTmp[16][8] , \u_div/CryTmp[16][7] ,
         \u_div/CryTmp[16][6] , \u_div/CryTmp[16][5] , \u_div/CryTmp[16][4] ,
         \u_div/CryTmp[16][3] , \u_div/CryTmp[16][2] , \u_div/CryTmp[16][23] ,
         \u_div/CryTmp[16][22] , \u_div/CryTmp[16][21] ,
         \u_div/CryTmp[16][20] , \u_div/CryTmp[16][19] ,
         \u_div/CryTmp[16][18] , \u_div/CryTmp[16][17] ,
         \u_div/CryTmp[16][16] , \u_div/CryTmp[16][15] ,
         \u_div/CryTmp[16][14] , \u_div/CryTmp[16][13] ,
         \u_div/CryTmp[16][12] , \u_div/CryTmp[16][11] ,
         \u_div/CryTmp[16][10] , \u_div/CryTmp[15][9] , \u_div/CryTmp[15][8] ,
         \u_div/CryTmp[15][7] , \u_div/CryTmp[15][6] , \u_div/CryTmp[15][5] ,
         \u_div/CryTmp[15][4] , \u_div/CryTmp[15][3] , \u_div/CryTmp[15][2] ,
         \u_div/CryTmp[15][24] , \u_div/CryTmp[15][23] ,
         \u_div/CryTmp[15][22] , \u_div/CryTmp[15][21] ,
         \u_div/CryTmp[15][20] , \u_div/CryTmp[15][19] ,
         \u_div/CryTmp[15][18] , \u_div/CryTmp[15][17] ,
         \u_div/CryTmp[15][16] , \u_div/CryTmp[15][15] ,
         \u_div/CryTmp[15][14] , \u_div/CryTmp[15][13] ,
         \u_div/CryTmp[15][12] , \u_div/CryTmp[15][11] ,
         \u_div/CryTmp[15][10] , net52402, net52401, net38340, net31107,
         net31046, net30917, net30665, net30662, net30607,
         \u_div/SumTmp[20][23] , \u_div/SumTmp[19][23] ,
         \u_div/SumTmp[19][22] , \u_div/SumTmp[19][21] ,
         \u_div/SumTmp[19][20] , \u_div/SumTmp[19][19] ,
         \u_div/SumTmp[19][18] , \u_div/SumTmp[19][16] ,
         \u_div/SumTmp[18][23] , \u_div/SumTmp[18][22] ,
         \u_div/SumTmp[18][21] , \u_div/SumTmp[18][20] ,
         \u_div/SumTmp[18][19] , \u_div/SumTmp[18][18] ,
         \u_div/SumTmp[18][17] , \u_div/SumTmp[17][23] ,
         \u_div/SumTmp[17][22] , \u_div/SumTmp[17][21] ,
         \u_div/SumTmp[17][20] , \u_div/SumTmp[17][0] ,
         \u_div/PartRem[21][23] , \u_div/PartRem[21][22] ,
         \u_div/PartRem[21][21] , \u_div/PartRem[21][20] ,
         \u_div/PartRem[21][19] , \u_div/PartRem[21][18] ,
         \u_div/PartRem[21][17] , \u_div/PartRem[20][24] ,
         \u_div/PartRem[20][23] , \u_div/PartRem[20][22] ,
         \u_div/PartRem[20][21] , \u_div/PartRem[20][20] ,
         \u_div/PartRem[20][19] , \u_div/PartRem[20][18] ,
         \u_div/PartRem[19][9] , \u_div/PartRem[19][8] ,
         \u_div/PartRem[19][7] , \u_div/PartRem[19][6] ,
         \u_div/PartRem[19][5] , \u_div/PartRem[19][4] ,
         \u_div/PartRem[19][3] , \u_div/PartRem[19][2] ,
         \u_div/PartRem[19][24] , \u_div/PartRem[19][23] ,
         \u_div/PartRem[19][22] , \u_div/PartRem[19][21] ,
         \u_div/PartRem[19][20] , \u_div/PartRem[19][1] ,
         \u_div/PartRem[19][19] , \u_div/PartRem[19][18] ,
         \u_div/PartRem[19][16] , \u_div/PartRem[19][15] ,
         \u_div/PartRem[19][14] , \u_div/PartRem[19][13] ,
         \u_div/PartRem[19][12] , \u_div/PartRem[19][11] ,
         \u_div/PartRem[19][10] , \u_div/PartRem[18][9] ,
         \u_div/PartRem[18][8] , \u_div/PartRem[18][7] ,
         \u_div/PartRem[18][6] , \u_div/PartRem[18][5] ,
         \u_div/PartRem[18][4] , \u_div/PartRem[18][3] ,
         \u_div/PartRem[18][2] , \u_div/PartRem[18][24] ,
         \u_div/PartRem[18][22] , \u_div/PartRem[18][21] ,
         \u_div/PartRem[18][20] , \u_div/PartRem[18][1] ,
         \u_div/PartRem[18][19] , \u_div/PartRem[18][18] ,
         \u_div/PartRem[18][17] , \u_div/PartRem[18][16] ,
         \u_div/PartRem[18][15] , \u_div/PartRem[18][14] ,
         \u_div/PartRem[18][13] , \u_div/PartRem[18][12] ,
         \u_div/PartRem[18][11] , \u_div/PartRem[18][10] ,
         \u_div/PartRem[17][1] , \u_div/CryTmp[20][23] ,
         \u_div/CryTmp[20][22] , \u_div/CryTmp[20][21] ,
         \u_div/CryTmp[20][20] , \u_div/CryTmp[20][19] ,
         \u_div/CryTmp[20][18] , \u_div/CryTmp[19][24] ,
         \u_div/CryTmp[19][23] , \u_div/CryTmp[19][22] ,
         \u_div/CryTmp[19][21] , \u_div/CryTmp[19][20] ,
         \u_div/CryTmp[19][19] , \u_div/CryTmp[18][9] , \u_div/CryTmp[18][8] ,
         \u_div/CryTmp[18][7] , \u_div/CryTmp[18][6] , \u_div/CryTmp[18][5] ,
         \u_div/CryTmp[18][4] , \u_div/CryTmp[18][3] , \u_div/CryTmp[18][2] ,
         \u_div/CryTmp[18][24] , \u_div/CryTmp[18][23] ,
         \u_div/CryTmp[18][22] , \u_div/CryTmp[18][21] ,
         \u_div/CryTmp[18][20] , \u_div/CryTmp[18][19] ,
         \u_div/CryTmp[18][18] , \u_div/CryTmp[18][17] ,
         \u_div/CryTmp[18][16] , \u_div/CryTmp[18][15] ,
         \u_div/CryTmp[18][14] , \u_div/CryTmp[18][13] ,
         \u_div/CryTmp[18][12] , \u_div/CryTmp[18][11] ,
         \u_div/CryTmp[18][10] , \u_div/CryTmp[17][9] , \u_div/CryTmp[17][8] ,
         \u_div/CryTmp[17][7] , \u_div/CryTmp[17][6] , \u_div/CryTmp[17][5] ,
         \u_div/CryTmp[17][4] , \u_div/CryTmp[17][3] , \u_div/CryTmp[17][2] ,
         \u_div/CryTmp[17][24] , \u_div/CryTmp[17][23] ,
         \u_div/CryTmp[17][22] , \u_div/CryTmp[17][21] ,
         \u_div/CryTmp[17][20] , \u_div/CryTmp[17][19] ,
         \u_div/CryTmp[17][18] , \u_div/CryTmp[17][17] ,
         \u_div/CryTmp[17][16] , \u_div/CryTmp[17][15] ,
         \u_div/CryTmp[17][14] , \u_div/CryTmp[17][13] ,
         \u_div/CryTmp[17][12] , \u_div/CryTmp[17][11] ,
         \u_div/CryTmp[17][10] , net38346, net38344, net30918, net30823,
         net30727, net30725, net30561, net30517, net30283, net30282, net30281,
         net30280, net30279, net30278, net30277, net30275, net30273, net30244,
         net30243, net30242, net30241, net30240, net30239, net30238, net30237,
         net30229, \*cell*33699/net34155 , \u_div/SumTmp[24][21] ,
         \u_div/SumTmp[24][20] , \u_div/SumTmp[23][23] ,
         \u_div/SumTmp[23][22] , \u_div/SumTmp[22][5] , \u_div/SumTmp[22][4] ,
         \u_div/SumTmp[21][9] , \u_div/SumTmp[21][8] , \u_div/SumTmp[21][7] ,
         \u_div/SumTmp[21][6] , \u_div/SumTmp[21][11] , \u_div/SumTmp[21][10] ,
         \u_div/SumTmp[20][16] , \u_div/SumTmp[20][15] ,
         \u_div/SumTmp[20][14] , \u_div/SumTmp[20][13] ,
         \u_div/SumTmp[20][12] , \u_div/SumTmp[19][17] ,
         \u_div/PartRem[25][21] , \u_div/PartRem[25][20] ,
         \u_div/PartRem[24][9] , \u_div/PartRem[24][8] ,
         \u_div/PartRem[24][7] , \u_div/PartRem[24][6] ,
         \u_div/PartRem[24][5] , \u_div/PartRem[24][4] ,
         \u_div/PartRem[24][3] , \u_div/PartRem[24][2] ,
         \u_div/PartRem[24][22] , \u_div/PartRem[24][21] ,
         \u_div/PartRem[24][20] , \u_div/PartRem[24][1] ,
         \u_div/PartRem[24][19] , \u_div/PartRem[24][18] ,
         \u_div/PartRem[24][17] , \u_div/PartRem[24][16] ,
         \u_div/PartRem[24][15] , \u_div/PartRem[24][14] ,
         \u_div/PartRem[24][13] , \u_div/PartRem[24][12] ,
         \u_div/PartRem[24][11] , \u_div/PartRem[24][10] ,
         \u_div/PartRem[23][5] , \u_div/PartRem[23][4] ,
         \u_div/PartRem[23][3] , \u_div/PartRem[23][2] ,
         \u_div/PartRem[23][24] , \u_div/PartRem[23][22] ,
         \u_div/PartRem[23][21] , \u_div/PartRem[23][20] ,
         \u_div/PartRem[23][1] , \u_div/PartRem[23][19] ,
         \u_div/PartRem[23][18] , \u_div/PartRem[23][17] ,
         \u_div/PartRem[22][9] , \u_div/PartRem[22][8] ,
         \u_div/PartRem[22][7] , \u_div/PartRem[22][6] ,
         \u_div/PartRem[22][4] , \u_div/PartRem[22][3] ,
         \u_div/PartRem[22][2] , \u_div/PartRem[22][1] ,
         \u_div/PartRem[22][11] , \u_div/PartRem[22][10] ,
         \u_div/PartRem[21][9] , \u_div/PartRem[21][7] ,
         \u_div/PartRem[21][6] , \u_div/PartRem[21][5] ,
         \u_div/PartRem[21][4] , \u_div/PartRem[21][3] ,
         \u_div/PartRem[21][2] , \u_div/PartRem[21][16] ,
         \u_div/PartRem[21][15] , \u_div/PartRem[21][14] ,
         \u_div/PartRem[21][13] , \u_div/PartRem[21][12] ,
         \u_div/PartRem[21][11] , \u_div/PartRem[21][10] ,
         \u_div/PartRem[20][9] , \u_div/PartRem[20][8] ,
         \u_div/PartRem[20][7] , \u_div/PartRem[20][6] ,
         \u_div/PartRem[20][5] , \u_div/PartRem[20][4] ,
         \u_div/PartRem[20][3] , \u_div/PartRem[20][2] ,
         \u_div/PartRem[20][1] , \u_div/PartRem[20][17] ,
         \u_div/PartRem[20][16] , \u_div/PartRem[20][15] ,
         \u_div/PartRem[20][14] , \u_div/PartRem[20][13] ,
         \u_div/PartRem[20][12] , \u_div/PartRem[20][11] ,
         \u_div/PartRem[20][10] , \u_div/CryTmp[24][22] ,
         \u_div/CryTmp[24][21] , \u_div/CryTmp[23][9] , \u_div/CryTmp[23][8] ,
         \u_div/CryTmp[23][7] , \u_div/CryTmp[23][6] , \u_div/CryTmp[23][5] ,
         \u_div/CryTmp[23][4] , \u_div/CryTmp[23][3] , \u_div/CryTmp[23][2] ,
         \u_div/CryTmp[23][23] , \u_div/CryTmp[23][22] ,
         \u_div/CryTmp[23][21] , \u_div/CryTmp[23][20] , \u_div/CryTmp[23][1] ,
         \u_div/CryTmp[23][19] , \u_div/CryTmp[23][18] ,
         \u_div/CryTmp[23][17] , \u_div/CryTmp[23][16] ,
         \u_div/CryTmp[23][15] , \u_div/CryTmp[23][14] ,
         \u_div/CryTmp[23][13] , \u_div/CryTmp[23][12] ,
         \u_div/CryTmp[23][11] , \u_div/CryTmp[23][10] , \u_div/CryTmp[22][5] ,
         \u_div/CryTmp[22][4] , \u_div/CryTmp[22][3] , \u_div/CryTmp[22][2] ,
         \u_div/CryTmp[22][24] , \u_div/CryTmp[22][23] ,
         \u_div/CryTmp[22][22] , \u_div/CryTmp[22][21] ,
         \u_div/CryTmp[22][20] , \u_div/CryTmp[22][19] ,
         \u_div/CryTmp[22][18] , \u_div/CryTmp[22][17] , \u_div/CryTmp[21][9] ,
         \u_div/CryTmp[21][8] , \u_div/CryTmp[21][7] , \u_div/CryTmp[21][6] ,
         \u_div/CryTmp[21][5] , \u_div/CryTmp[21][4] , \u_div/CryTmp[21][3] ,
         \u_div/CryTmp[21][2] , \u_div/CryTmp[21][12] , \u_div/CryTmp[21][11] ,
         \u_div/CryTmp[21][10] , \u_div/CryTmp[20][9] , \u_div/CryTmp[20][8] ,
         \u_div/CryTmp[20][7] , \u_div/CryTmp[20][6] , \u_div/CryTmp[20][5] ,
         \u_div/CryTmp[20][4] , \u_div/CryTmp[20][3] , \u_div/CryTmp[20][2] ,
         \u_div/CryTmp[20][17] , \u_div/CryTmp[20][16] ,
         \u_div/CryTmp[20][15] , \u_div/CryTmp[20][14] ,
         \u_div/CryTmp[20][13] , \u_div/CryTmp[20][12] ,
         \u_div/CryTmp[20][11] , \u_div/CryTmp[20][10] , \u_div/CryTmp[19][9] ,
         \u_div/CryTmp[19][8] , \u_div/CryTmp[19][7] , \u_div/CryTmp[19][6] ,
         \u_div/CryTmp[19][5] , \u_div/CryTmp[19][4] , \u_div/CryTmp[19][3] ,
         \u_div/CryTmp[19][2] , \u_div/CryTmp[19][18] , \u_div/CryTmp[19][17] ,
         \u_div/CryTmp[19][16] , \u_div/CryTmp[19][15] ,
         \u_div/CryTmp[19][14] , \u_div/CryTmp[19][13] ,
         \u_div/CryTmp[19][12] , \u_div/CryTmp[19][11] ,
         \u_div/CryTmp[19][10] , n1240, net31094, net31074, net31052, net31030,
         net31007, net30983, net30982, net30956, net30872, net30824, net30776,
         net30775, net30201, net30189, net30188, net30179, net30138, net30137,
         net30136, net30134, net30133, net30132, net30131, net30045, net30044,
         net30041, net30040, net30039, net30038, net30037, net30035, net30032,
         net30031, net30030, net30029, net30028, net30027, net30026, net30025,
         \u_div/SumTmp[26][8] , \u_div/SumTmp[25][9] , \u_div/SumTmp[25][21] ,
         \u_div/SumTmp[25][20] , \u_div/SumTmp[25][19] ,
         \u_div/SumTmp[25][18] , \u_div/SumTmp[25][17] ,
         \u_div/SumTmp[25][16] , \u_div/SumTmp[25][15] ,
         \u_div/SumTmp[25][14] , \u_div/SumTmp[25][13] ,
         \u_div/SumTmp[25][12] , \u_div/SumTmp[25][11] ,
         \u_div/SumTmp[25][10] , \u_div/SumTmp[24][19] ,
         \u_div/SumTmp[24][18] , \u_div/SumTmp[24][17] ,
         \u_div/SumTmp[24][16] , \u_div/SumTmp[24][15] ,
         \u_div/SumTmp[24][14] , \u_div/PartRem[26][9] ,
         \u_div/PartRem[26][8] , \u_div/PartRem[26][7] ,
         \u_div/PartRem[26][6] , \u_div/PartRem[26][5] ,
         \u_div/PartRem[26][4] , \u_div/PartRem[26][3] ,
         \u_div/PartRem[26][2] , \u_div/PartRem[26][21] ,
         \u_div/PartRem[26][20] , \u_div/PartRem[26][1] ,
         \u_div/PartRem[26][19] , \u_div/PartRem[26][18] ,
         \u_div/PartRem[26][17] , \u_div/PartRem[26][16] ,
         \u_div/PartRem[26][15] , \u_div/PartRem[26][14] ,
         \u_div/PartRem[26][13] , \u_div/PartRem[26][12] ,
         \u_div/PartRem[26][11] , \u_div/PartRem[26][10] ,
         \u_div/PartRem[25][9] , \u_div/PartRem[25][8] ,
         \u_div/PartRem[25][7] , \u_div/PartRem[25][6] ,
         \u_div/PartRem[25][5] , \u_div/PartRem[25][4] ,
         \u_div/PartRem[25][3] , \u_div/PartRem[25][2] ,
         \u_div/PartRem[25][19] , \u_div/PartRem[25][18] ,
         \u_div/PartRem[25][17] , \u_div/PartRem[25][16] ,
         \u_div/PartRem[25][15] , \u_div/PartRem[25][14] ,
         \u_div/PartRem[25][13] , \u_div/PartRem[25][12] ,
         \u_div/PartRem[25][11] , \u_div/PartRem[25][10] ,
         \u_div/CryTmp[25][9] , \u_div/CryTmp[25][8] , \u_div/CryTmp[25][7] ,
         \u_div/CryTmp[25][6] , \u_div/CryTmp[25][5] , \u_div/CryTmp[25][4] ,
         \u_div/CryTmp[25][3] , \u_div/CryTmp[25][2] , \u_div/CryTmp[25][22] ,
         \u_div/CryTmp[25][21] , \u_div/CryTmp[25][20] , \u_div/CryTmp[25][1] ,
         \u_div/CryTmp[25][19] , \u_div/CryTmp[25][18] ,
         \u_div/CryTmp[25][17] , \u_div/CryTmp[25][16] ,
         \u_div/CryTmp[25][15] , \u_div/CryTmp[25][14] ,
         \u_div/CryTmp[25][13] , \u_div/CryTmp[25][12] ,
         \u_div/CryTmp[25][11] , \u_div/CryTmp[25][10] , \u_div/CryTmp[24][9] ,
         \u_div/CryTmp[24][8] , \u_div/CryTmp[24][7] , \u_div/CryTmp[24][6] ,
         \u_div/CryTmp[24][5] , \u_div/CryTmp[24][4] , \u_div/CryTmp[24][3] ,
         \u_div/CryTmp[24][2] , \u_div/CryTmp[24][20] , \u_div/CryTmp[24][1] ,
         \u_div/CryTmp[24][19] , \u_div/CryTmp[24][18] ,
         \u_div/CryTmp[24][17] , \u_div/CryTmp[24][16] ,
         \u_div/CryTmp[24][15] , \u_div/CryTmp[24][14] ,
         \u_div/CryTmp[24][13] , \u_div/CryTmp[24][12] ,
         \u_div/CryTmp[24][11] , \u_div/CryTmp[24][10] , net31317, net31315,
         net30878, net30877, net30829, net30781, net30685, net30684, net30637,
         net30589, net30541, net30493, net30250, net30024, net30023, net30021,
         net30020, net30019, net30018, net30017, net30016, net30014, net30011,
         net30010, net30009, net30008, net30007, net30006, net30005, net30004,
         net30003, net30001, net30000, net29999, net29998, net29997, net29996,
         net29995, net29994, net29993, net29992, net29991, net29990, net29989,
         net29988, net29987, net29986, net29985, net29984,
         \u_div/SumTmp[29][17] , \u_div/SumTmp[28][9] , \u_div/SumTmp[28][8] ,
         \u_div/SumTmp[28][7] , \u_div/SumTmp[28][6] , \u_div/SumTmp[28][5] ,
         \u_div/SumTmp[28][4] , \u_div/SumTmp[28][3] , \u_div/SumTmp[28][2] ,
         \u_div/SumTmp[28][1] , \u_div/SumTmp[27][10] , \u_div/SumTmp[26][20] ,
         \u_div/SumTmp[26][19] , \u_div/SumTmp[26][18] ,
         \u_div/SumTmp[26][17] , \u_div/SumTmp[26][16] ,
         \u_div/SumTmp[26][15] , \u_div/SumTmp[26][14] ,
         \u_div/SumTmp[26][13] , \u_div/SumTmp[26][12] ,
         \u_div/SumTmp[26][11] , \u_div/PartRem[30][9] ,
         \u_div/PartRem[30][8] , \u_div/PartRem[30][7] ,
         \u_div/PartRem[30][6] , \u_div/PartRem[30][5] ,
         \u_div/PartRem[30][4] , \u_div/PartRem[30][3] ,
         \u_div/PartRem[30][2] , \u_div/PartRem[30][1] ,
         \u_div/PartRem[30][17] , \u_div/PartRem[30][16] ,
         \u_div/PartRem[30][15] , \u_div/PartRem[30][14] ,
         \u_div/PartRem[30][13] , \u_div/PartRem[30][12] ,
         \u_div/PartRem[30][11] , \u_div/PartRem[30][10] ,
         \u_div/PartRem[29][9] , \u_div/PartRem[29][8] ,
         \u_div/PartRem[29][7] , \u_div/PartRem[29][6] ,
         \u_div/PartRem[29][5] , \u_div/PartRem[29][4] ,
         \u_div/PartRem[29][3] , \u_div/PartRem[29][2] ,
         \u_div/PartRem[29][1] , \u_div/PartRem[28][9] ,
         \u_div/PartRem[28][8] , \u_div/PartRem[28][7] ,
         \u_div/PartRem[28][6] , \u_div/PartRem[28][5] ,
         \u_div/PartRem[28][4] , \u_div/PartRem[28][3] ,
         \u_div/PartRem[28][2] , \u_div/PartRem[28][1] ,
         \u_div/PartRem[28][10] , \u_div/PartRem[27][9] ,
         \u_div/PartRem[27][8] , \u_div/PartRem[27][7] ,
         \u_div/PartRem[27][6] , \u_div/PartRem[27][5] ,
         \u_div/PartRem[27][4] , \u_div/PartRem[27][3] ,
         \u_div/PartRem[27][2] , \u_div/PartRem[27][20] ,
         \u_div/PartRem[27][1] , \u_div/PartRem[27][19] ,
         \u_div/PartRem[27][18] , \u_div/PartRem[27][17] ,
         \u_div/PartRem[27][16] , \u_div/PartRem[27][15] ,
         \u_div/PartRem[27][14] , \u_div/PartRem[27][13] ,
         \u_div/PartRem[27][12] , \u_div/PartRem[27][11] ,
         \u_div/PartRem[27][10] , \u_div/CryTmp[29][9] , \u_div/CryTmp[29][8] ,
         \u_div/CryTmp[29][7] , \u_div/CryTmp[29][6] , \u_div/CryTmp[29][5] ,
         \u_div/CryTmp[29][4] , \u_div/CryTmp[29][3] , \u_div/CryTmp[29][2] ,
         \u_div/CryTmp[29][1] , \u_div/CryTmp[29][18] , \u_div/CryTmp[29][17] ,
         \u_div/CryTmp[29][16] , \u_div/CryTmp[29][15] ,
         \u_div/CryTmp[29][14] , \u_div/CryTmp[29][13] ,
         \u_div/CryTmp[29][12] , \u_div/CryTmp[29][11] ,
         \u_div/CryTmp[29][10] , \u_div/CryTmp[28][9] , \u_div/CryTmp[28][8] ,
         \u_div/CryTmp[28][7] , \u_div/CryTmp[28][6] , \u_div/CryTmp[28][5] ,
         \u_div/CryTmp[28][4] , \u_div/CryTmp[28][3] , \u_div/CryTmp[28][2] ,
         \u_div/CryTmp[28][1] , \u_div/CryTmp[28][10] , \u_div/CryTmp[27][9] ,
         \u_div/CryTmp[27][8] , \u_div/CryTmp[27][7] , \u_div/CryTmp[27][6] ,
         \u_div/CryTmp[27][5] , \u_div/CryTmp[27][4] , \u_div/CryTmp[27][3] ,
         \u_div/CryTmp[27][2] , \u_div/CryTmp[27][1] , \u_div/CryTmp[27][10] ,
         \u_div/CryTmp[26][9] , \u_div/CryTmp[26][8] , \u_div/CryTmp[26][7] ,
         \u_div/CryTmp[26][6] , \u_div/CryTmp[26][5] , \u_div/CryTmp[26][4] ,
         \u_div/CryTmp[26][3] , \u_div/CryTmp[26][2] , \u_div/CryTmp[26][21] ,
         \u_div/CryTmp[26][20] , \u_div/CryTmp[26][1] , \u_div/CryTmp[26][19] ,
         \u_div/CryTmp[26][18] , \u_div/CryTmp[26][17] ,
         \u_div/CryTmp[26][16] , \u_div/CryTmp[26][15] ,
         \u_div/CryTmp[26][14] , \u_div/CryTmp[26][13] ,
         \u_div/CryTmp[26][12] , \u_div/CryTmp[26][11] ,
         \u_div/CryTmp[26][10] , net49672, net30735, net30734, net30002,
         net29983, net29973, net29972, net29971, net29970, net29969, net29968,
         net29967, net29966, net29965, net29930, net29920, net29919, net29918,
         net29917, net29916, net29913, net29912, net29911, net29910, net29909,
         net29908, net29907, net29906, net29905, \u_div/SumTmp[36][3] ,
         \u_div/SumTmp[35][4] , \u_div/SumTmp[34][9] , \u_div/SumTmp[34][8] ,
         \u_div/SumTmp[34][7] , \u_div/SumTmp[34][6] , \u_div/SumTmp[34][5] ,
         \u_div/SumTmp[33][10] , \u_div/SumTmp[32][14] ,
         \u_div/SumTmp[32][13] , \u_div/SumTmp[32][12] ,
         \u_div/SumTmp[32][11] , \u_div/SumTmp[31][14] ,
         \u_div/SumTmp[30][16] , \u_div/SumTmp[30][15] ,
         \u_div/PartRem[37][3] , \u_div/PartRem[37][2] ,
         \u_div/PartRem[37][1] , \u_div/PartRem[36][4] ,
         \u_div/PartRem[36][2] , \u_div/PartRem[36][1] ,
         \u_div/PartRem[35][9] , \u_div/PartRem[35][7] ,
         \u_div/PartRem[35][6] , \u_div/PartRem[35][5] ,
         \u_div/PartRem[35][4] , \u_div/PartRem[35][3] ,
         \u_div/PartRem[35][2] , \u_div/PartRem[35][1] ,
         \u_div/PartRem[34][9] , \u_div/PartRem[34][8] ,
         \u_div/PartRem[34][7] , \u_div/PartRem[34][6] ,
         \u_div/PartRem[34][5] , \u_div/PartRem[34][4] ,
         \u_div/PartRem[34][3] , \u_div/PartRem[34][2] ,
         \u_div/PartRem[34][1] , \u_div/PartRem[34][10] ,
         \u_div/PartRem[33][9] , \u_div/PartRem[33][8] ,
         \u_div/PartRem[33][7] , \u_div/PartRem[33][6] ,
         \u_div/PartRem[33][5] , \u_div/PartRem[33][4] ,
         \u_div/PartRem[33][3] , \u_div/PartRem[33][2] ,
         \u_div/PartRem[33][1] , \u_div/PartRem[33][14] ,
         \u_div/PartRem[33][13] , \u_div/PartRem[33][12] ,
         \u_div/PartRem[33][11] , \u_div/PartRem[33][10] ,
         \u_div/PartRem[32][9] , \u_div/PartRem[32][8] ,
         \u_div/PartRem[32][7] , \u_div/PartRem[32][6] ,
         \u_div/PartRem[32][5] , \u_div/PartRem[32][4] ,
         \u_div/PartRem[32][3] , \u_div/PartRem[32][2] ,
         \u_div/PartRem[32][1] , \u_div/PartRem[32][14] ,
         \u_div/PartRem[32][13] , \u_div/PartRem[32][12] ,
         \u_div/PartRem[32][11] , \u_div/PartRem[32][10] ,
         \u_div/PartRem[31][9] , \u_div/PartRem[31][8] ,
         \u_div/PartRem[31][7] , \u_div/PartRem[31][6] ,
         \u_div/PartRem[31][5] , \u_div/PartRem[31][4] ,
         \u_div/PartRem[31][3] , \u_div/PartRem[31][2] ,
         \u_div/PartRem[31][1] , \u_div/PartRem[31][16] ,
         \u_div/PartRem[31][15] , \u_div/PartRem[31][14] ,
         \u_div/PartRem[31][13] , \u_div/PartRem[31][12] ,
         \u_div/PartRem[31][11] , \u_div/PartRem[31][10] ,
         \u_div/CryTmp[36][3] , \u_div/CryTmp[36][2] , \u_div/CryTmp[36][1] ,
         \u_div/CryTmp[35][4] , \u_div/CryTmp[35][3] , \u_div/CryTmp[35][2] ,
         \u_div/CryTmp[35][1] , \u_div/CryTmp[34][9] , \u_div/CryTmp[34][8] ,
         \u_div/CryTmp[34][7] , \u_div/CryTmp[34][6] , \u_div/CryTmp[34][5] ,
         \u_div/CryTmp[34][4] , \u_div/CryTmp[34][3] , \u_div/CryTmp[34][2] ,
         \u_div/CryTmp[34][1] , \u_div/CryTmp[34][10] , \u_div/CryTmp[33][9] ,
         \u_div/CryTmp[33][8] , \u_div/CryTmp[33][7] , \u_div/CryTmp[33][6] ,
         \u_div/CryTmp[33][5] , \u_div/CryTmp[33][4] , \u_div/CryTmp[33][3] ,
         \u_div/CryTmp[33][2] , \u_div/CryTmp[33][1] , \u_div/CryTmp[33][10] ,
         \u_div/CryTmp[32][9] , \u_div/CryTmp[32][8] , \u_div/CryTmp[32][7] ,
         \u_div/CryTmp[32][6] , \u_div/CryTmp[32][5] , \u_div/CryTmp[32][4] ,
         \u_div/CryTmp[32][3] , \u_div/CryTmp[32][2] , \u_div/CryTmp[32][1] ,
         \u_div/CryTmp[32][15] , \u_div/CryTmp[32][14] ,
         \u_div/CryTmp[32][13] , \u_div/CryTmp[32][12] ,
         \u_div/CryTmp[32][11] , \u_div/CryTmp[32][10] , \u_div/CryTmp[31][9] ,
         \u_div/CryTmp[31][8] , \u_div/CryTmp[31][7] , \u_div/CryTmp[31][6] ,
         \u_div/CryTmp[31][5] , \u_div/CryTmp[31][4] , \u_div/CryTmp[31][3] ,
         \u_div/CryTmp[31][2] , \u_div/CryTmp[31][1] , \u_div/CryTmp[31][14] ,
         \u_div/CryTmp[31][13] , \u_div/CryTmp[31][12] ,
         \u_div/CryTmp[31][11] , \u_div/CryTmp[31][10] , \u_div/CryTmp[30][9] ,
         \u_div/CryTmp[30][8] , \u_div/CryTmp[30][7] , \u_div/CryTmp[30][6] ,
         \u_div/CryTmp[30][5] , \u_div/CryTmp[30][4] , \u_div/CryTmp[30][3] ,
         \u_div/CryTmp[30][2] , \u_div/CryTmp[30][1] , \u_div/CryTmp[30][17] ,
         \u_div/CryTmp[30][16] , \u_div/CryTmp[30][15] ,
         \u_div/CryTmp[30][14] , \u_div/CryTmp[30][13] ,
         \u_div/CryTmp[30][12] , \u_div/CryTmp[30][11] ,
         \u_div/CryTmp[30][10] , net52311, net46015, net30148, net30147,
         net29904, net29903, net29902, net29901, net29900, net29898, net29897,
         net29896, net29895, net29894, net29893, net29892, net29891, net29890,
         net29836, net29828, \u_div/SumTmp[43][3] , \u_div/SumTmp[43][2] ,
         \u_div/SumTmp[43][1] , \u_div/SumTmp[42][4] , \u_div/SumTmp[41][5] ,
         \u_div/SumTmp[40][6] , \u_div/SumTmp[39][7] , \u_div/SumTmp[39][6] ,
         \u_div/SumTmp[38][8] , \u_div/SumTmp[38][7] , \u_div/SumTmp[38][1] ,
         \u_div/SumTmp[37][2] , \u_div/SumTmp[37][1] , \u_div/PartRem[45][2] ,
         \u_div/PartRem[45][1] , \u_div/PartRem[44][3] ,
         \u_div/PartRem[44][2] , \u_div/PartRem[44][1] ,
         \u_div/PartRem[43][4] , \u_div/PartRem[43][3] ,
         \u_div/PartRem[43][2] , \u_div/PartRem[43][1] ,
         \u_div/PartRem[42][5] , \u_div/PartRem[42][4] ,
         \u_div/PartRem[42][3] , \u_div/PartRem[42][2] ,
         \u_div/PartRem[41][6] , \u_div/PartRem[41][5] ,
         \u_div/PartRem[41][4] , \u_div/PartRem[41][3] ,
         \u_div/PartRem[41][2] , \u_div/PartRem[41][1] ,
         \u_div/PartRem[40][7] , \u_div/PartRem[40][6] ,
         \u_div/PartRem[40][5] , \u_div/PartRem[40][4] ,
         \u_div/PartRem[40][3] , \u_div/PartRem[40][2] ,
         \u_div/PartRem[40][1] , \u_div/PartRem[39][8] ,
         \u_div/PartRem[39][7] , \u_div/PartRem[39][4] ,
         \u_div/PartRem[39][3] , \u_div/PartRem[39][1] ,
         \u_div/PartRem[38][1] , \u_div/CryTmp[44][3] , \u_div/CryTmp[44][2] ,
         \u_div/CryTmp[44][1] , \u_div/CryTmp[43][4] , \u_div/CryTmp[43][3] ,
         \u_div/CryTmp[43][2] , \u_div/CryTmp[43][1] , \u_div/CryTmp[42][4] ,
         \u_div/CryTmp[42][3] , \u_div/CryTmp[42][2] , \u_div/CryTmp[42][1] ,
         \u_div/CryTmp[41][5] , \u_div/CryTmp[41][4] , \u_div/CryTmp[41][3] ,
         \u_div/CryTmp[41][2] , \u_div/CryTmp[41][1] , \u_div/CryTmp[40][6] ,
         \u_div/CryTmp[40][5] , \u_div/CryTmp[40][4] , \u_div/CryTmp[40][3] ,
         \u_div/CryTmp[40][2] , \u_div/CryTmp[40][1] , \u_div/CryTmp[39][8] ,
         \u_div/CryTmp[39][7] , \u_div/CryTmp[39][6] , \u_div/CryTmp[39][5] ,
         \u_div/CryTmp[39][4] , \u_div/CryTmp[39][3] , \u_div/CryTmp[39][2] ,
         \u_div/CryTmp[39][1] , \u_div/CryTmp[38][9] , \u_div/CryTmp[38][8] ,
         \u_div/CryTmp[38][7] , \u_div/CryTmp[38][6] , \u_div/CryTmp[38][5] ,
         \u_div/CryTmp[38][4] , \u_div/CryTmp[38][3] , \u_div/CryTmp[38][2] ,
         \u_div/CryTmp[38][1] , \u_div/CryTmp[37][3] , \u_div/CryTmp[37][2] ,
         \u_div/CryTmp[37][1] , net37262, net31546, net30697, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n174,
         n175, n176, n177, n178, n179, n180, n181, n182, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n985, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239;
  assign quotient[7] = net32518;
  assign quotient[10] = net32538;
  assign quotient[11] = net32544;
  assign quotient[17] = net32580;
  assign quotient[19] = net32590;
  assign quotient[20] = net32598;
  assign quotient[22] = net32610;
  assign quotient[37] = net37242;
  assign quotient[34] = net37563;
  assign quotient[36] = net37570;
  assign quotient[30] = net37577;
  assign quotient[38] = net37581;
  assign quotient[41] = net37584;
  assign quotient[33] = net37854;
  assign quotient[31] = net40084;
  assign quotient[6] = net40656;
  assign quotient[8] = net40719;
  assign quotient[27] = net41415;
  assign quotient[4] = net42040;
  assign quotient[13] = net42408;
  assign quotient[42] = net43819;
  assign quotient[3] = net45597;
  assign quotient[18] = net45665;
  assign quotient[9] = net46550;
  assign quotient[29] = net47679;
  assign quotient[24] = net47709;
  assign quotient[14] = net47718;
  assign quotient[32] = net50049;
  assign quotient[40] = net50182;
  assign quotient[35] = net50471;

  FADDX1_RVT \u_div/u_fa_PartRem_0_2_23  ( .A(net31800), .B(
        \u_div/CryTmp[2][23] ), .CI(\u_div/PartRem[3][23] ), .CO(
        \u_div/CryTmp[2][24] ), .S(\u_div/SumTmp[2][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_19  ( .A(\u_div/PartRem[2][19] ), .B(
        net31910), .CI(\u_div/CryTmp[1][19] ), .CO(\u_div/CryTmp[1][20] ), .S(
        \u_div/SumTmp[1][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_23  ( .A(n908), .B(net31800), .CI(n220), 
        .CO(\u_div/CryTmp[0][24] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_19  ( .A(\u_div/PartRem[1][19] ), .B(
        net31910), .CI(n942), .CO(\u_div/CryTmp[0][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_11  ( .A(\u_div/PartRem[35][11] ), .B(
        net49055), .CI(net44064), .CO(\u_div/CryTmp[34][12] ), .S(
        \u_div/SumTmp[34][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_21  ( .A(\u_div/PartRem[1][21] ), .B(
        net31854), .CI(n926), .CO(\u_div/CryTmp[0][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_22  ( .A(n910), .B(net31826), .CI(n922), 
        .CO(\u_div/CryTmp[0][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_15  ( .A(n972), .B(net32012), .CI(n977), 
        .CO(\u_div/CryTmp[0][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_16  ( .A(n970), .B(net31986), .CI(
        \u_div/CryTmp[0][16] ), .CO(\u_div/CryTmp[0][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_12  ( .A(\u_div/PartRem[28][12] ), .B(
        net32088), .CI(\u_div/CryTmp[27][12] ), .CO(\u_div/CryTmp[27][13] ), 
        .S(\u_div/SumTmp[27][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_13  ( .A(net49679), .B(net32078), .CI(
        n906), .CO(\u_div/CryTmp[27][14] ), .S(\u_div/SumTmp[27][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_15  ( .A(\u_div/PartRem[29][15] ), .B(
        net32016), .CI(\u_div/CryTmp[28][15] ), .CO(\u_div/CryTmp[28][16] ), 
        .S(\u_div/SumTmp[28][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_11  ( .A(\u_div/PartRem[28][11] ), .B(
        net49055), .CI(\u_div/CryTmp[27][11] ), .CO(\u_div/CryTmp[27][12] ), 
        .S(\u_div/SumTmp[27][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_21  ( .A(\u_div/PartRem[3][21] ), .B(
        net31854), .CI(\u_div/CryTmp[2][21] ), .CO(\u_div/CryTmp[2][22] ), .S(
        \u_div/SumTmp[2][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_11  ( .A(\u_div/PartRem[34][11] ), .B(
        net49055), .CI(\u_div/CryTmp[33][11] ), .CO(\u_div/CryTmp[33][12] ), 
        .S(\u_div/SumTmp[33][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_6  ( .A(\u_div/PartRem[38][6] ), .B(
        net32272), .CI(\u_div/CryTmp[37][6] ), .CO(\u_div/CryTmp[37][7] ), .S(
        \u_div/SumTmp[37][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_4  ( .A(\u_div/PartRem[38][4] ), .B(
        net32326), .CI(\u_div/CryTmp[37][4] ), .CO(\u_div/CryTmp[37][5] ), .S(
        \u_div/SumTmp[37][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_5  ( .A(\u_div/PartRem[38][5] ), .B(
        net32302), .CI(\u_div/CryTmp[37][5] ), .CO(\u_div/CryTmp[37][6] ), .S(
        \u_div/SumTmp[37][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_8  ( .A(\u_div/PartRem[37][8] ), .B(
        net32196), .CI(\u_div/CryTmp[36][8] ), .CO(\u_div/CryTmp[36][9] ), .S(
        \u_div/SumTmp[36][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_7  ( .A(\u_div/PartRem[36][7] ), .B(
        net32242), .CI(\u_div/CryTmp[35][7] ), .CO(\u_div/CryTmp[35][8] ), .S(
        \u_div/SumTmp[35][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_4  ( .A(\u_div/PartRem[37][4] ), .B(
        net32326), .CI(\u_div/CryTmp[36][4] ), .CO(\u_div/CryTmp[36][5] ), .S(
        \u_div/SumTmp[36][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_5  ( .A(\u_div/PartRem[37][5] ), .B(
        net32302), .CI(\u_div/CryTmp[36][5] ), .CO(\u_div/CryTmp[36][6] ), .S(
        \u_div/SumTmp[36][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_17  ( .A(n966), .B(net31964), .CI(n272), 
        .CO(\u_div/CryTmp[0][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_13  ( .A(\u_div/PartRem[1][13] ), .B(
        net32068), .CI(\u_div/CryTmp[0][13] ), .CO(\u_div/CryTmp[0][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_14  ( .A(\u_div/PartRem[1][14] ), .B(
        net32042), .CI(\u_div/CryTmp[0][14] ), .CO(\u_div/CryTmp[0][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_11  ( .A(\u_div/PartRem[29][11] ), .B(
        net49055), .CI(\u_div/CryTmp[28][11] ), .CO(\u_div/CryTmp[28][12] ), 
        .S(\u_div/SumTmp[28][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_10  ( .A(\u_div/PartRem[29][10] ), .B(
        net32140), .CI(net42939), .CO(\u_div/CryTmp[28][11] ), .S(
        \u_div/SumTmp[28][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_6  ( .A(\u_div/PartRem[36][6] ), .B(
        net32254), .CI(n1001), .CO(\u_div/CryTmp[35][7] ), .S(
        \u_div/SumTmp[35][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_11  ( .A(\u_div/PartRem[1][11] ), .B(
        net32118), .CI(\u_div/CryTmp[0][11] ), .CO(\u_div/CryTmp[0][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_12  ( .A(\u_div/PartRem[1][12] ), .B(
        net32092), .CI(\u_div/CryTmp[0][12] ), .CO(\u_div/CryTmp[0][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_3  ( .A(n274), .B(net32354), .CI(
        net46242), .CO(\u_div/CryTmp[37][4] ), .S(\u_div/SumTmp[37][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_1  ( .A(\u_div/PartRem[1][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[0][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_2  ( .A(\u_div/PartRem[1][2] ), .B(
        net32362), .CI(\u_div/CryTmp[0][2] ), .CO(\u_div/CryTmp[0][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_3  ( .A(\u_div/PartRem[1][3] ), .B(
        net32334), .CI(\u_div/CryTmp[0][3] ), .CO(\u_div/CryTmp[0][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_1  ( .A(\u_div/PartRem[2][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[1][2] ), .S(
        \u_div/SumTmp[1][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_1  ( .A(\u_div/PartRem[3][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[2][2] ), .S(
        \u_div/SumTmp[2][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_8  ( .A(\u_div/PartRem[1][8] ), .B(
        net32196), .CI(\u_div/CryTmp[0][8] ), .CO(\u_div/CryTmp[0][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_9  ( .A(\u_div/PartRem[1][9] ), .B(
        net32168), .CI(\u_div/CryTmp[0][9] ), .CO(\u_div/CryTmp[0][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_4  ( .A(\u_div/PartRem[1][4] ), .B(
        net32310), .CI(\u_div/CryTmp[0][4] ), .CO(\u_div/CryTmp[0][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_5  ( .A(\u_div/PartRem[1][5] ), .B(
        net32280), .CI(\u_div/CryTmp[0][5] ), .CO(\u_div/CryTmp[0][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_10  ( .A(\u_div/PartRem[1][10] ), .B(
        net32144), .CI(\u_div/CryTmp[0][10] ), .CO(\u_div/CryTmp[0][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_13  ( .A(\u_div/PartRem[29][13] ), .B(
        net32078), .CI(n107), .CO(\u_div/CryTmp[28][14] ), .S(
        \u_div/SumTmp[28][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_17  ( .A(\u_div/PartRem[29][17] ), .B(
        net31960), .CI(n892), .CO(\u_div/CryTmp[28][18] ), .S(
        \u_div/SumTmp[28][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_10  ( .A(\u_div/PartRem[2][10] ), .B(
        net32144), .CI(\u_div/CryTmp[1][10] ), .CO(\u_div/CryTmp[1][11] ), .S(
        \u_div/SumTmp[1][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_2  ( .A(\u_div/PartRem[2][2] ), .B(
        net32362), .CI(\u_div/CryTmp[1][2] ), .CO(\u_div/CryTmp[1][3] ), .S(
        \u_div/SumTmp[1][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_4  ( .A(\u_div/PartRem[2][4] ), .B(
        net32310), .CI(\u_div/CryTmp[1][4] ), .CO(\u_div/CryTmp[1][5] ), .S(
        \u_div/SumTmp[1][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_11  ( .A(n982), .B(net32118), .CI(
        \u_div/CryTmp[1][11] ), .CO(\u_div/CryTmp[1][12] ), .S(
        \u_div/SumTmp[1][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_14  ( .A(\u_div/PartRem[2][14] ), .B(
        net32042), .CI(n924), .CO(\u_div/CryTmp[1][15] ), .S(
        \u_div/SumTmp[1][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_18  ( .A(\u_div/PartRem[2][18] ), .B(
        net31938), .CI(\u_div/CryTmp[1][18] ), .CO(\u_div/CryTmp[1][19] ), .S(
        \u_div/SumTmp[1][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_14  ( .A(\u_div/PartRem[29][14] ), .B(
        net32046), .CI(\u_div/CryTmp[28][14] ), .CO(\u_div/CryTmp[28][15] ), 
        .S(\u_div/SumTmp[28][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_11  ( .A(\u_div/PartRem[7][11] ), .B(
        net32118), .CI(\u_div/CryTmp[6][11] ), .CO(\u_div/CryTmp[6][12] ), .S(
        \u_div/SumTmp[6][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_10  ( .A(\u_div/PartRem[7][10] ), .B(
        net32144), .CI(net49281), .CO(\u_div/CryTmp[6][11] ), .S(
        \u_div/SumTmp[6][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_11  ( .A(n1003), .B(net32118), .CI(
        \u_div/CryTmp[7][11] ), .CO(\u_div/CryTmp[7][12] ), .S(
        \u_div/SumTmp[7][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_10  ( .A(\u_div/PartRem[8][10] ), .B(
        net32144), .CI(\u_div/CryTmp[7][10] ), .CO(\u_div/CryTmp[7][11] ), .S(
        \u_div/SumTmp[7][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_11  ( .A(\u_div/PartRem[23][11] ), .B(
        net32116), .CI(\u_div/CryTmp[22][11] ), .CO(\u_div/CryTmp[22][12] ), 
        .S(\u_div/SumTmp[22][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_10  ( .A(\u_div/PartRem[23][10] ), .B(
        net32142), .CI(\u_div/CryTmp[22][10] ), .CO(\u_div/CryTmp[22][11] ), 
        .S(\u_div/SumTmp[22][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_8  ( .A(\u_div/PartRem[23][8] ), .B(
        net32198), .CI(\u_div/CryTmp[22][8] ), .CO(\u_div/CryTmp[22][9] ), .S(
        \u_div/SumTmp[22][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_13  ( .A(\u_div/PartRem[3][13] ), .B(
        net32068), .CI(\u_div/CryTmp[2][13] ), .CO(\u_div/CryTmp[2][14] ), .S(
        \u_div/SumTmp[2][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_14  ( .A(\u_div/PartRem[3][14] ), .B(
        net32042), .CI(\u_div/CryTmp[2][14] ), .CO(\u_div/CryTmp[2][15] ), .S(
        \u_div/SumTmp[2][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_17  ( .A(\u_div/PartRem[3][17] ), .B(
        net31964), .CI(\u_div/CryTmp[2][17] ), .CO(\u_div/CryTmp[2][18] ), .S(
        \u_div/SumTmp[2][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_18  ( .A(\u_div/PartRem[3][18] ), .B(
        net31940), .CI(\u_div/CryTmp[2][18] ), .CO(\u_div/CryTmp[2][19] ), .S(
        \u_div/SumTmp[2][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_13  ( .A(\u_div/PartRem[23][13] ), .B(
        net32066), .CI(\u_div/CryTmp[22][13] ), .CO(\u_div/CryTmp[22][14] ), 
        .S(\u_div/SumTmp[22][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_13  ( .A(\u_div/PartRem[7][13] ), .B(
        net32068), .CI(\u_div/CryTmp[6][13] ), .CO(\u_div/CryTmp[6][14] ), .S(
        \u_div/SumTmp[6][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_8  ( .A(\u_div/PartRem[38][8] ), .B(
        net32212), .CI(n940), .CO(\u_div/CryTmp[37][9] ), .S(
        \u_div/SumTmp[37][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_13  ( .A(\u_div/PartRem[8][13] ), .B(
        net32068), .CI(\u_div/CryTmp[7][13] ), .CO(\u_div/CryTmp[7][14] ), .S(
        \u_div/SumTmp[7][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_14  ( .A(\u_div/PartRem[7][14] ), .B(
        net32042), .CI(\u_div/CryTmp[6][14] ), .CO(\u_div/CryTmp[6][15] ), .S(
        \u_div/SumTmp[6][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_17  ( .A(\u_div/PartRem[22][17] ), .B(
        net31960), .CI(\u_div/CryTmp[21][17] ), .CO(\u_div/CryTmp[21][18] ), 
        .S(\u_div/SumTmp[21][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_10  ( .A(\u_div/PartRem[3][10] ), .B(
        net32144), .CI(\u_div/CryTmp[2][10] ), .CO(\u_div/CryTmp[2][11] ), .S(
        \u_div/SumTmp[2][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_14  ( .A(\u_div/PartRem[28][14] ), .B(
        net32046), .CI(\u_div/CryTmp[27][14] ), .CO(\u_div/CryTmp[27][15] ), 
        .S(\u_div/SumTmp[27][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_17  ( .A(n324), .B(net31960), .CI(
        \u_div/CryTmp[27][17] ), .CO(\u_div/CryTmp[27][18] ), .S(
        \u_div/SumTmp[27][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_14  ( .A(\u_div/PartRem[22][14] ), .B(
        net32044), .CI(\u_div/CryTmp[21][14] ), .CO(\u_div/CryTmp[21][15] ), 
        .S(\u_div/SumTmp[21][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_14  ( .A(\u_div/PartRem[8][14] ), .B(
        net32042), .CI(\u_div/CryTmp[7][14] ), .CO(\u_div/CryTmp[7][15] ), .S(
        \u_div/SumTmp[7][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_2  ( .A(\u_div/PartRem[3][2] ), .B(
        net32362), .CI(\u_div/CryTmp[2][2] ), .CO(\u_div/CryTmp[2][3] ), .S(
        \u_div/SumTmp[2][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_4  ( .A(\u_div/PartRem[3][4] ), .B(
        net32310), .CI(\u_div/CryTmp[2][4] ), .CO(\u_div/CryTmp[2][5] ), .S(
        \u_div/SumTmp[2][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_8  ( .A(n936), .B(net32196), .CI(n957), 
        .CO(\u_div/CryTmp[2][9] ), .S(\u_div/SumTmp[2][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_13  ( .A(n40), .B(net32078), .CI(n932), 
        .CO(\u_div/CryTmp[33][14] ), .S(\u_div/SumTmp[33][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_10  ( .A(\u_div/PartRem[37][10] ), .B(
        net32140), .CI(\u_div/CryTmp[36][10] ), .CO(\u_div/CryTmp[36][11] ), 
        .S(\u_div/SumTmp[36][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_22  ( .A(\u_div/PartRem[25][22] ), .B(
        net31826), .CI(net48534), .CO(\u_div/CryTmp[24][23] ), .S(
        \u_div/SumTmp[24][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_6  ( .A(\u_div/PartRem[1][6] ), .B(
        net32250), .CI(\u_div/CryTmp[0][6] ), .CO(\u_div/CryTmp[0][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_7  ( .A(\u_div/PartRem[1][7] ), .B(
        net32226), .CI(\u_div/CryTmp[0][7] ), .CO(\u_div/CryTmp[0][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_3  ( .A(\u_div/PartRem[2][3] ), .B(
        net32334), .CI(\u_div/CryTmp[1][3] ), .CO(\u_div/CryTmp[1][4] ), .S(
        \u_div/SumTmp[1][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_5  ( .A(\u_div/PartRem[2][5] ), .B(
        net32280), .CI(\u_div/CryTmp[1][5] ), .CO(\u_div/CryTmp[1][6] ), .S(
        \u_div/SumTmp[1][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_6  ( .A(\u_div/PartRem[2][6] ), .B(
        net32250), .CI(\u_div/CryTmp[1][6] ), .CO(\u_div/CryTmp[1][7] ), .S(
        \u_div/SumTmp[1][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_7  ( .A(\u_div/PartRem[2][7] ), .B(
        net32226), .CI(\u_div/CryTmp[1][7] ), .CO(\u_div/CryTmp[1][8] ), .S(
        \u_div/SumTmp[1][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_9  ( .A(\u_div/PartRem[2][9] ), .B(
        net32168), .CI(n955), .CO(\u_div/CryTmp[1][10] ), .S(
        \u_div/SumTmp[1][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_20  ( .A(\u_div/PartRem[2][20] ), .B(
        net31882), .CI(\u_div/CryTmp[1][20] ), .CO(\u_div/CryTmp[1][21] ), .S(
        \u_div/SumTmp[1][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_15  ( .A(\u_div/PartRem[2][15] ), .B(
        net32012), .CI(\u_div/CryTmp[1][15] ), .CO(\u_div/CryTmp[1][16] ), .S(
        \u_div/SumTmp[1][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_16  ( .A(\u_div/PartRem[2][16] ), .B(
        net31986), .CI(n222), .CO(\u_div/CryTmp[1][17] ), .S(
        \u_div/SumTmp[1][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_12  ( .A(n1010), .B(\u_div/CryTmp[1][12] ), .CI(net32092), .CO(\u_div/CryTmp[1][13] ), .S(\u_div/SumTmp[1][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_12  ( .A(\u_div/PartRem[3][12] ), .B(n918), .CI(net32092), .CO(\u_div/CryTmp[2][13] ), .S(\u_div/SumTmp[2][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_7  ( .A(\u_div/PartRem[37][7] ), .B(
        net32242), .CI(n992), .CO(\u_div/CryTmp[36][8] ), .S(
        \u_div/SumTmp[36][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_12  ( .A(n38), .B(n42), .CI(net32092), 
        .CO(\u_div/CryTmp[6][13] ), .S(\u_div/SumTmp[6][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_12  ( .A(\u_div/PartRem[8][12] ), .B(
        net32092), .CI(n266), .CO(\u_div/CryTmp[7][13] ), .S(
        \u_div/SumTmp[7][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_9  ( .A(\u_div/PartRem[8][9] ), .B(
        net32168), .CI(\u_div/CryTmp[7][9] ), .CO(\u_div/CryTmp[7][10] ), .S(
        \u_div/SumTmp[7][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_12  ( .A(\u_div/PartRem[23][12] ), .B(
        net32090), .CI(\u_div/CryTmp[22][12] ), .CO(\u_div/CryTmp[22][13] ), 
        .S(\u_div/SumTmp[22][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_9  ( .A(\u_div/PartRem[23][9] ), .B(
        net32166), .CI(\u_div/CryTmp[22][9] ), .CO(\u_div/CryTmp[22][10] ), 
        .S(\u_div/SumTmp[22][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_7  ( .A(\u_div/PartRem[23][7] ), .B(
        net32222), .CI(\u_div/CryTmp[22][7] ), .CO(\u_div/CryTmp[22][8] ), .S(
        \u_div/SumTmp[22][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_6  ( .A(\u_div/PartRem[23][6] ), .B(
        net32252), .CI(\u_div/CryTmp[22][6] ), .CO(\u_div/CryTmp[22][7] ), .S(
        \u_div/SumTmp[22][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_9  ( .A(\u_div/PartRem[3][9] ), .B(
        net32168), .CI(\u_div/CryTmp[2][9] ), .CO(\u_div/CryTmp[2][10] ), .S(
        \u_div/SumTmp[2][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_15  ( .A(\u_div/PartRem[3][15] ), .B(
        net32012), .CI(\u_div/CryTmp[2][15] ), .CO(\u_div/CryTmp[2][16] ), .S(
        \u_div/SumTmp[2][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_16  ( .A(\u_div/PartRem[3][16] ), .B(
        net31986), .CI(n920), .CO(\u_div/CryTmp[2][17] ), .S(
        \u_div/SumTmp[2][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_21  ( .A(\u_div/PartRem[22][21] ), .B(
        net31856), .CI(n228), .CO(\u_div/CryTmp[21][22] ), .S(
        \u_div/SumTmp[21][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_15  ( .A(\u_div/PartRem[28][15] ), .B(
        net32016), .CI(\u_div/CryTmp[27][15] ), .CO(\u_div/CryTmp[27][16] ), 
        .S(\u_div/SumTmp[27][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_16  ( .A(\u_div/PartRem[28][16] ), .B(
        net31982), .CI(\u_div/CryTmp[27][16] ), .CO(\u_div/CryTmp[27][17] ), 
        .S(\u_div/SumTmp[27][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_12  ( .A(n71), .B(net32090), .CI(
        net49113), .CO(\u_div/CryTmp[21][13] ), .S(\u_div/SumTmp[21][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_21  ( .A(\u_div/PartRem[15][21] ), .B(
        net31856), .CI(net48639), .CO(\u_div/CryTmp[14][22] ), .S(
        \u_div/SumTmp[14][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_21  ( .A(\u_div/PartRem[14][21] ), .B(
        net31856), .CI(\u_div/CryTmp[13][21] ), .CO(\u_div/CryTmp[13][22] ), 
        .S(\u_div/SumTmp[13][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_15  ( .A(\u_div/PartRem[7][15] ), .B(
        net32012), .CI(\u_div/CryTmp[6][15] ), .CO(\u_div/CryTmp[6][16] ), .S(
        \u_div/SumTmp[6][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_15  ( .A(\u_div/PartRem[8][15] ), .B(
        net32012), .CI(\u_div/CryTmp[7][15] ), .CO(\u_div/CryTmp[7][16] ), .S(
        \u_div/SumTmp[7][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_16  ( .A(\u_div/PartRem[7][16] ), .B(
        net31986), .CI(\u_div/CryTmp[6][16] ), .CO(\u_div/CryTmp[6][17] ), .S(
        \u_div/SumTmp[6][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_16  ( .A(\u_div/PartRem[8][16] ), .B(
        net31984), .CI(n944), .CO(\u_div/CryTmp[7][17] ), .S(
        \u_div/SumTmp[7][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_19  ( .A(\u_div/PartRem[7][19] ), .B(
        net31910), .CI(\u_div/CryTmp[6][19] ), .CO(\u_div/CryTmp[6][20] ), .S(
        \u_div/SumTmp[6][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_21  ( .A(\u_div/PartRem[7][21] ), .B(
        net31854), .CI(n930), .CO(\u_div/CryTmp[6][22] ), .S(
        \u_div/SumTmp[6][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_3  ( .A(\u_div/PartRem[3][3] ), .B(
        net32334), .CI(\u_div/CryTmp[2][3] ), .CO(\u_div/CryTmp[2][4] ), .S(
        \u_div/SumTmp[2][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_5  ( .A(\u_div/PartRem[3][5] ), .B(
        net32280), .CI(\u_div/CryTmp[2][5] ), .CO(\u_div/CryTmp[2][6] ), .S(
        \u_div/SumTmp[2][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_6  ( .A(\u_div/PartRem[3][6] ), .B(
        net32250), .CI(n997), .CO(\u_div/CryTmp[2][7] ), .S(
        \u_div/SumTmp[2][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_7  ( .A(\u_div/PartRem[3][7] ), .B(
        net32226), .CI(\u_div/CryTmp[2][7] ), .CO(\u_div/CryTmp[2][8] ), .S(
        \u_div/SumTmp[2][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_19  ( .A(\u_div/PartRem[3][19] ), .B(
        net31910), .CI(n902), .CO(\u_div/CryTmp[2][20] ), .S(
        \u_div/SumTmp[2][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_20  ( .A(\u_div/PartRem[3][20] ), .B(
        net31882), .CI(\u_div/CryTmp[2][20] ), .CO(\u_div/CryTmp[2][21] ), .S(
        \u_div/SumTmp[2][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_19  ( .A(net44395), .B(n994), .CI(
        net31914), .CO(\u_div/CryTmp[27][20] ), .S(\u_div/SumTmp[27][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_9  ( .A(\u_div/PartRem[38][9] ), .B(
        net32186), .CI(\u_div/CryTmp[37][9] ), .CO(\u_div/CryTmp[37][10] ), 
        .S(\u_div/SumTmp[37][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_15  ( .A(\u_div/PartRem[22][15] ), .B(
        net32014), .CI(n270), .CO(\u_div/CryTmp[21][16] ), .S(
        \u_div/SumTmp[21][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_23  ( .A(n1009), .B(net31800), .CI(
        \u_div/CryTmp[5][23] ), .CO(\u_div/CryTmp[5][24] ), .S(
        \u_div/SumTmp[5][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_23  ( .A(\u_div/PartRem[7][23] ), .B(
        net31800), .CI(\u_div/CryTmp[6][23] ), .CO(\u_div/CryTmp[6][24] ), .S(
        \u_div/SumTmp[6][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_23  ( .A(\u_div/PartRem[10][23] ), .B(
        net31800), .CI(n968), .CO(\u_div/CryTmp[9][24] ), .S(
        \u_div/SumTmp[9][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_23  ( .A(\u_div/PartRem[14][23] ), .B(
        net31802), .CI(n127), .CO(\u_div/CryTmp[13][24] ), .S(
        \u_div/SumTmp[13][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_23  ( .A(\u_div/PartRem[15][23] ), .B(
        net31802), .CI(\u_div/CryTmp[14][23] ), .CO(\u_div/CryTmp[14][24] ), 
        .S(\u_div/SumTmp[14][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_18  ( .A(\u_div/PartRem[7][18] ), .B(
        net31940), .CI(n885), .CO(\u_div/CryTmp[6][19] ), .S(
        \u_div/SumTmp[6][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_18  ( .A(\u_div/PartRem[22][18] ), .B(
        net31938), .CI(\u_div/CryTmp[21][18] ), .CO(\u_div/CryTmp[21][19] ), 
        .S(\u_div/SumTmp[21][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_22  ( .A(\u_div/PartRem[7][22] ), .B(
        net31826), .CI(\u_div/CryTmp[6][22] ), .CO(\u_div/CryTmp[6][23] ), .S(
        \u_div/SumTmp[6][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_22  ( .A(\u_div/PartRem[22][22] ), .B(
        net31828), .CI(\u_div/CryTmp[21][22] ), .CO(\u_div/CryTmp[21][23] ), 
        .S(\u_div/SumTmp[21][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_20  ( .A(\u_div/PartRem[10][20] ), .B(
        net31882), .CI(\u_div/CryTmp[9][20] ), .CO(\u_div/CryTmp[9][21] ), .S(
        \u_div/SumTmp[9][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_20  ( .A(\u_div/PartRem[7][20] ), .B(
        net31882), .CI(\u_div/CryTmp[6][20] ), .CO(\u_div/CryTmp[6][21] ), .S(
        \u_div/SumTmp[6][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_22  ( .A(\u_div/PartRem[15][22] ), .B(
        net31828), .CI(\u_div/CryTmp[14][22] ), .CO(\u_div/CryTmp[14][23] ), 
        .S(\u_div/SumTmp[14][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_22  ( .A(\u_div/PartRem[10][22] ), .B(
        net31826), .CI(\u_div/CryTmp[9][22] ), .CO(\u_div/CryTmp[9][23] ), .S(
        \u_div/SumTmp[9][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_20  ( .A(\u_div/PartRem[22][20] ), .B(
        net31884), .CI(n1005), .CO(\u_div/CryTmp[21][21] ), .S(
        \u_div/SumTmp[21][20] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_21_19  ( .A(\u_div/PartRem[22][19] ), .B(
        net31912), .CI(n900), .CO(\u_div/CryTmp[21][20] ), .S(
        \u_div/SumTmp[21][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_18  ( .A(\u_div/PartRem[29][18] ), .B(
        net31940), .CI(n990), .CO(\u_div/CryTmp[28][19] ), .S(
        \u_div/SumTmp[28][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_18  ( .A(\u_div/PartRem[28][18] ), .B(
        net31938), .CI(\u_div/CryTmp[27][18] ), .CO(\u_div/CryTmp[27][19] ), 
        .S(\u_div/SumTmp[27][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_23  ( .A(\u_div/PartRem[22][23] ), .B(
        net31802), .CI(\u_div/CryTmp[21][23] ), .CO(\u_div/CryTmp[21][24] ), 
        .S(\u_div/SumTmp[21][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_11  ( .A(n1011), .B(net32118), .CI(
        \u_div/CryTmp[2][11] ), .CO(\u_div/CryTmp[2][12] ), .S(
        \u_div/SumTmp[2][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_2_22  ( .A(\u_div/PartRem[3][22] ), .B(
        net31826), .CI(\u_div/CryTmp[2][22] ), .CO(\u_div/CryTmp[2][23] ), .S(
        \u_div/SumTmp[2][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_16  ( .A(\u_div/PartRem[22][16] ), .B(
        net31982), .CI(n69), .CO(\u_div/CryTmp[21][17] ), .S(
        \u_div/SumTmp[21][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_9  ( .A(\u_div/PartRem[36][9] ), .B(
        net32186), .CI(n928), .CO(\u_div/CryTmp[35][10] ), .S(
        \u_div/SumTmp[35][9] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_37_7  ( .A(\u_div/PartRem[38][7] ), .B(
        net32226), .CI(\u_div/CryTmp[37][7] ), .CO(\u_div/CryTmp[37][8] ), .S(
        \u_div/SumTmp[37][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_8  ( .A(\u_div/PartRem[36][8] ), .B(
        net32200), .CI(\u_div/CryTmp[35][8] ), .CO(\u_div/CryTmp[35][9] ), .S(
        \u_div/SumTmp[35][8] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_31_15  ( .A(\u_div/PartRem[32][15] ), .B(
        net32016), .CI(net42398), .CO(\u_div/CryTmp[31][16] ), .S(
        \u_div/SumTmp[31][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_17  ( .A(\u_div/PartRem[8][17] ), .B(
        net31962), .CI(n262), .CO(\u_div/CryTmp[7][18] ), .S(
        \u_div/SumTmp[7][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_19  ( .A(\u_div/PartRem[8][19] ), .B(
        net31910), .CI(\u_div/CryTmp[7][19] ), .CO(\u_div/CryTmp[7][20] ), .S(
        \u_div/SumTmp[7][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_21  ( .A(n855), .B(net31854), .CI(
        \u_div/CryTmp[7][21] ), .CO(\u_div/CryTmp[7][22] ), .S(
        \u_div/SumTmp[7][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_22  ( .A(\u_div/PartRem[8][22] ), .B(
        net31826), .CI(\u_div/CryTmp[7][22] ), .CO(\u_div/CryTmp[7][23] ), .S(
        \u_div/SumTmp[7][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_23  ( .A(\u_div/PartRem[8][23] ), .B(
        net31800), .CI(\u_div/CryTmp[7][23] ), .CO(\u_div/CryTmp[7][24] ), .S(
        \u_div/SumTmp[7][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_20  ( .A(\u_div/PartRem[9][20] ), .B(
        net31882), .CI(\u_div/CryTmp[8][20] ), .CO(\u_div/CryTmp[8][21] ), .S(
        \u_div/SumTmp[8][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_21  ( .A(\u_div/PartRem[9][21] ), .B(
        net31854), .CI(\u_div/CryTmp[8][21] ), .CO(\u_div/CryTmp[8][22] ), .S(
        \u_div/SumTmp[8][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_22  ( .A(\u_div/PartRem[9][22] ), .B(
        net31826), .CI(\u_div/CryTmp[8][22] ), .CO(\u_div/CryTmp[8][23] ), .S(
        \u_div/SumTmp[8][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_23  ( .A(\u_div/PartRem[9][23] ), .B(
        net31800), .CI(\u_div/CryTmp[8][23] ), .CO(\u_div/CryTmp[8][24] ), .S(
        \u_div/SumTmp[8][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_1  ( .A(net32382), .B(
        \u_div/PartRem[8][1] ), .CI(\u_div/CryTmp[11][1] ), .CO(
        \u_div/CryTmp[7][2] ), .S(\u_div/SumTmp[7][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_2  ( .A(\u_div/PartRem[8][2] ), .B(
        net32362), .CI(\u_div/CryTmp[7][2] ), .CO(\u_div/CryTmp[7][3] ), .S(
        \u_div/SumTmp[7][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_3  ( .A(\u_div/PartRem[8][3] ), .B(
        net32334), .CI(\u_div/CryTmp[7][3] ), .CO(\u_div/CryTmp[7][4] ), .S(
        \u_div/SumTmp[7][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_4  ( .A(\u_div/PartRem[8][4] ), .B(
        net32310), .CI(\u_div/CryTmp[7][4] ), .CO(\u_div/CryTmp[7][5] ), .S(
        \u_div/SumTmp[7][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_5  ( .A(\u_div/PartRem[8][5] ), .B(
        net32280), .CI(\u_div/CryTmp[7][5] ), .CO(\u_div/CryTmp[7][6] ), .S(
        \u_div/SumTmp[7][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_6  ( .A(\u_div/PartRem[8][6] ), .B(
        net32250), .CI(\u_div/CryTmp[7][6] ), .CO(\u_div/CryTmp[7][7] ), .S(
        \u_div/SumTmp[7][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_7  ( .A(net40783), .B(net32224), .CI(
        \u_div/CryTmp[7][7] ), .CO(\u_div/CryTmp[7][8] ), .S(
        \u_div/SumTmp[7][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_8  ( .A(\u_div/PartRem[8][8] ), .B(
        net32196), .CI(n264), .CO(\u_div/CryTmp[7][9] ), .S(
        \u_div/SumTmp[7][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_1  ( .A(\u_div/PartRem[7][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[6][2] ), .S(
        \u_div/SumTmp[6][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_2  ( .A(\u_div/PartRem[7][2] ), .B(
        net32362), .CI(\u_div/CryTmp[6][2] ), .CO(\u_div/CryTmp[6][3] ), .S(
        \u_div/SumTmp[6][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_3  ( .A(\u_div/PartRem[7][3] ), .B(
        net32334), .CI(\u_div/CryTmp[6][3] ), .CO(\u_div/CryTmp[6][4] ), .S(
        \u_div/SumTmp[6][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_4  ( .A(n880), .B(net32310), .CI(n878), 
        .CO(\u_div/CryTmp[6][5] ), .S(\u_div/SumTmp[6][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_5  ( .A(n882), .B(net32280), .CI(
        \u_div/CryTmp[6][5] ), .CO(\u_div/CryTmp[6][6] ), .S(
        \u_div/SumTmp[6][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_6  ( .A(n853), .B(net32250), .CI(
        \u_div/PartRem[7][6] ), .CO(\u_div/CryTmp[6][7] ), .S(
        \u_div/SumTmp[6][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_7  ( .A(\u_div/PartRem[7][7] ), .B(
        net32224), .CI(\u_div/CryTmp[6][7] ), .CO(\u_div/CryTmp[6][8] ), .S(
        \u_div/SumTmp[6][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_8  ( .A(\u_div/PartRem[7][8] ), .B(
        net32196), .CI(\u_div/CryTmp[6][8] ), .CO(\u_div/CryTmp[6][9] ), .S(
        \u_div/SumTmp[6][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_9  ( .A(\u_div/PartRem[7][9] ), .B(
        net32168), .CI(\u_div/CryTmp[6][9] ), .CO(\u_div/CryTmp[6][10] ), .S(
        \u_div/SumTmp[6][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_22  ( .A(net38272), .B(net31826), .CI(
        n216), .CO(\u_div/CryTmp[5][23] ), .S(\u_div/SumTmp[5][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_1  ( .A(\u_div/PartRem[6][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[5][2] ), .S(
        \u_div/SumTmp[5][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_2  ( .A(\u_div/PartRem[6][2] ), .B(
        net32362), .CI(\u_div/CryTmp[5][2] ), .CO(\u_div/CryTmp[5][3] ), .S(
        \u_div/SumTmp[5][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_3  ( .A(\u_div/PartRem[6][3] ), .B(
        net32334), .CI(\u_div/CryTmp[5][3] ), .CO(\u_div/CryTmp[5][4] ), .S(
        \u_div/SumTmp[5][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_4  ( .A(\u_div/PartRem[6][4] ), .B(
        net32310), .CI(\u_div/CryTmp[5][4] ), .CO(\u_div/CryTmp[5][5] ), .S(
        \u_div/SumTmp[5][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_5  ( .A(\u_div/PartRem[6][5] ), .B(
        net32280), .CI(n849), .CO(\u_div/CryTmp[5][6] ), .S(
        \u_div/SumTmp[5][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_6  ( .A(\u_div/PartRem[6][6] ), .B(
        net32250), .CI(n851), .CO(\u_div/CryTmp[5][7] ), .S(
        \u_div/SumTmp[5][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_7  ( .A(\u_div/CryTmp[5][7] ), .B(
        net32224), .CI(n874), .CO(\u_div/CryTmp[5][8] ), .S(
        \u_div/SumTmp[5][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_8  ( .A(net52000), .B(net32196), .CI(
        \u_div/CryTmp[5][8] ), .CO(\u_div/CryTmp[5][9] ), .S(
        \u_div/SumTmp[5][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_9  ( .A(net52003), .B(net32168), .CI(
        \u_div/CryTmp[5][9] ), .CO(\u_div/CryTmp[5][10] ), .S(
        \u_div/SumTmp[5][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_10  ( .A(n875), .B(net32144), .CI(
        \u_div/CryTmp[5][10] ), .CO(\u_div/CryTmp[5][11] ), .S(
        \u_div/SumTmp[5][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_11  ( .A(\u_div/PartRem[6][11] ), .B(
        net32118), .CI(\u_div/CryTmp[5][11] ), .CO(\u_div/CryTmp[5][12] ), .S(
        \u_div/SumTmp[5][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_12  ( .A(\u_div/PartRem[6][12] ), .B(
        \u_div/CryTmp[5][12] ), .CI(net32092), .CO(\u_div/CryTmp[5][13] ), .S(
        \u_div/SumTmp[5][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_13  ( .A(\u_div/PartRem[6][13] ), .B(
        net32068), .CI(\u_div/CryTmp[5][13] ), .CO(\u_div/CryTmp[5][14] ), .S(
        \u_div/SumTmp[5][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_14  ( .A(\u_div/PartRem[6][14] ), .B(
        net32042), .CI(\u_div/CryTmp[5][14] ), .CO(\u_div/CryTmp[5][15] ), .S(
        \u_div/SumTmp[5][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_15  ( .A(\u_div/PartRem[6][15] ), .B(
        net32012), .CI(n89), .CO(\u_div/CryTmp[5][16] ), .S(
        \u_div/SumTmp[5][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_16  ( .A(\u_div/PartRem[6][16] ), .B(
        net31986), .CI(\u_div/CryTmp[5][16] ), .CO(\u_div/CryTmp[5][17] ), .S(
        \u_div/SumTmp[5][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_17  ( .A(\u_div/PartRem[6][17] ), .B(
        net31964), .CI(\u_div/CryTmp[5][17] ), .CO(\u_div/CryTmp[5][18] ), .S(
        \u_div/SumTmp[5][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_18  ( .A(\u_div/PartRem[6][18] ), .B(
        net31940), .CI(\u_div/CryTmp[5][18] ), .CO(\u_div/CryTmp[5][19] ), .S(
        \u_div/SumTmp[5][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_19  ( .A(\u_div/PartRem[6][19] ), .B(
        net31910), .CI(\u_div/CryTmp[5][19] ), .CO(\u_div/CryTmp[5][20] ), .S(
        \u_div/SumTmp[5][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_5_20  ( .A(\u_div/PartRem[6][20] ), .B(
        net31882), .CI(\u_div/CryTmp[5][20] ), .CO(\u_div/CryTmp[5][21] ), .S(
        \u_div/SumTmp[5][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_1  ( .A(\u_div/PartRem[5][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[4][2] ), .S(
        \u_div/SumTmp[4][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_2  ( .A(\u_div/PartRem[5][2] ), .B(
        net32362), .CI(\u_div/CryTmp[4][2] ), .CO(\u_div/CryTmp[4][3] ), .S(
        \u_div/SumTmp[4][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_3  ( .A(\u_div/PartRem[5][3] ), .B(
        net32334), .CI(\u_div/CryTmp[4][3] ), .CO(\u_div/CryTmp[4][4] ), .S(
        \u_div/SumTmp[4][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_5  ( .A(\u_div/PartRem[5][5] ), .B(
        net32280), .CI(n841), .CO(\u_div/CryTmp[4][6] ), .S(
        \u_div/SumTmp[4][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_6  ( .A(\u_div/PartRem[5][6] ), .B(
        net32250), .CI(n252), .CO(\u_div/CryTmp[4][7] ), .S(
        \u_div/SumTmp[4][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_7  ( .A(n869), .B(net32224), .CI(n868), 
        .CO(\u_div/CryTmp[4][8] ), .S(\u_div/SumTmp[4][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_8  ( .A(\u_div/PartRem[5][8] ), .B(
        net32196), .CI(\u_div/CryTmp[4][8] ), .CO(\u_div/CryTmp[4][9] ), .S(
        \u_div/SumTmp[4][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_9  ( .A(\u_div/PartRem[5][9] ), .B(
        net32168), .CI(\u_div/CryTmp[4][9] ), .CO(\u_div/CryTmp[4][10] ), .S(
        \u_div/SumTmp[4][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_10  ( .A(\u_div/PartRem[5][10] ), .B(
        net32144), .CI(\u_div/CryTmp[4][10] ), .CO(\u_div/CryTmp[4][11] ), .S(
        \u_div/SumTmp[4][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_12  ( .A(\u_div/PartRem[5][12] ), .B(
        net32092), .CI(n67), .CO(\u_div/CryTmp[4][13] ), .S(
        \u_div/SumTmp[4][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_13  ( .A(\u_div/PartRem[5][13] ), .B(
        net32068), .CI(\u_div/CryTmp[4][13] ), .CO(\u_div/CryTmp[4][14] ), .S(
        \u_div/SumTmp[4][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_14  ( .A(\u_div/PartRem[5][14] ), .B(
        net32042), .CI(\u_div/CryTmp[4][14] ), .CO(\u_div/CryTmp[4][15] ), .S(
        \u_div/SumTmp[4][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_15  ( .A(\u_div/PartRem[5][15] ), .B(
        net32012), .CI(\u_div/CryTmp[4][15] ), .CO(\u_div/CryTmp[4][16] ), .S(
        \u_div/SumTmp[4][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_16  ( .A(\u_div/PartRem[5][16] ), .B(
        net31986), .CI(\u_div/CryTmp[4][16] ), .CO(\u_div/CryTmp[4][17] ), .S(
        \u_div/SumTmp[4][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_17  ( .A(\u_div/PartRem[5][17] ), .B(
        net31964), .CI(\u_div/CryTmp[4][17] ), .CO(\u_div/CryTmp[4][18] ), .S(
        \u_div/SumTmp[4][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_19  ( .A(n125), .B(net31910), .CI(n268), 
        .CO(\u_div/CryTmp[4][20] ), .S(\u_div/SumTmp[4][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_20  ( .A(\u_div/PartRem[5][20] ), .B(
        net31882), .CI(n870), .CO(\u_div/CryTmp[4][21] ), .S(
        \u_div/SumTmp[4][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_21  ( .A(\u_div/PartRem[5][21] ), .B(
        net31854), .CI(n859), .CO(\u_div/CryTmp[4][22] ), .S(
        \u_div/SumTmp[4][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_22  ( .A(n873), .B(net31826), .CI(
        \u_div/CryTmp[4][22] ), .CO(\u_div/CryTmp[4][23] ), .S(
        \u_div/SumTmp[4][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_23  ( .A(n836), .B(net31800), .CI(n77), 
        .CO(\u_div/CryTmp[4][24] ), .S(\u_div/SumTmp[4][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_1  ( .A(\u_div/PartRem[4][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[3][2] ), .S(
        \u_div/SumTmp[3][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_2  ( .A(\u_div/PartRem[4][2] ), .B(
        net32362), .CI(n276), .CO(\u_div/CryTmp[3][3] ), .S(
        \u_div/SumTmp[3][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_3  ( .A(\u_div/PartRem[4][3] ), .B(
        net32334), .CI(\u_div/CryTmp[3][3] ), .CO(\u_div/CryTmp[3][4] ), .S(
        \u_div/SumTmp[3][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_4  ( .A(\u_div/PartRem[4][4] ), .B(
        net32310), .CI(n258), .CO(\u_div/CryTmp[3][5] ), .S(
        \u_div/SumTmp[3][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_6  ( .A(n844), .B(net32250), .CI(
        \u_div/PartRem[4][6] ), .CO(\u_div/CryTmp[3][7] ), .S(
        \u_div/SumTmp[3][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_7  ( .A(\u_div/PartRem[4][7] ), .B(
        net32226), .CI(\u_div/CryTmp[3][7] ), .CO(\u_div/CryTmp[3][8] ), .S(
        \u_div/SumTmp[3][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_8  ( .A(\u_div/PartRem[4][8] ), .B(
        net32196), .CI(n846), .CO(\u_div/CryTmp[3][9] ), .S(
        \u_div/SumTmp[3][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_9  ( .A(\u_div/PartRem[4][9] ), .B(
        net32168), .CI(\u_div/CryTmp[3][9] ), .CO(\u_div/CryTmp[3][10] ), .S(
        \u_div/SumTmp[3][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_10  ( .A(\u_div/PartRem[4][10] ), .B(
        net32144), .CI(n861), .CO(\u_div/CryTmp[3][11] ), .S(
        \u_div/SumTmp[3][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_13  ( .A(\u_div/PartRem[4][13] ), .B(
        net32068), .CI(\u_div/CryTmp[3][13] ), .CO(\u_div/CryTmp[3][14] ), .S(
        \u_div/SumTmp[3][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_14  ( .A(\u_div/PartRem[4][14] ), .B(
        net32042), .CI(n865), .CO(\u_div/CryTmp[3][15] ), .S(
        \u_div/SumTmp[3][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_15  ( .A(\u_div/PartRem[4][15] ), .B(
        net32012), .CI(\u_div/CryTmp[3][15] ), .CO(\u_div/CryTmp[3][16] ), .S(
        \u_div/SumTmp[3][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_16  ( .A(\u_div/PartRem[4][16] ), .B(
        net31986), .CI(\u_div/CryTmp[3][16] ), .CO(\u_div/CryTmp[3][17] ), .S(
        \u_div/SumTmp[3][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_17  ( .A(\u_div/PartRem[4][17] ), .B(
        net31964), .CI(\u_div/CryTmp[3][17] ), .CO(\u_div/CryTmp[3][18] ), .S(
        \u_div/SumTmp[3][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_18  ( .A(\u_div/PartRem[4][18] ), .B(
        net31938), .CI(\u_div/CryTmp[3][18] ), .CO(\u_div/CryTmp[3][19] ), .S(
        \u_div/SumTmp[3][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_20  ( .A(\u_div/PartRem[4][20] ), .B(
        net31882), .CI(\u_div/CryTmp[3][20] ), .CO(\u_div/CryTmp[3][21] ), .S(
        \u_div/SumTmp[3][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_22  ( .A(\u_div/PartRem[4][22] ), .B(
        net31826), .CI(\u_div/CryTmp[3][22] ), .CO(\u_div/CryTmp[3][23] ), .S(
        \u_div/SumTmp[3][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_23  ( .A(net31800), .B(n867), .CI(
        net50743), .CO(\u_div/CryTmp[3][24] ), .S(\u_div/SumTmp[3][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_17  ( .A(\u_div/PartRem[11][17] ), .B(
        net31962), .CI(\u_div/CryTmp[10][17] ), .CO(\u_div/CryTmp[10][18] ), 
        .S(\u_div/SumTmp[10][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_18  ( .A(\u_div/PartRem[11][18] ), .B(
        net31940), .CI(\u_div/CryTmp[10][18] ), .CO(\u_div/CryTmp[10][19] ), 
        .S(\u_div/SumTmp[10][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_20  ( .A(\u_div/PartRem[11][20] ), .B(
        n300), .CI(net31882), .CO(\u_div/CryTmp[10][21] ), .S(
        \u_div/SumTmp[10][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_21  ( .A(\u_div/PartRem[11][21] ), .B(
        net31854), .CI(n79), .CO(\u_div/CryTmp[10][22] ), .S(
        \u_div/SumTmp[10][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_22  ( .A(\u_div/PartRem[11][22] ), .B(
        net31826), .CI(\u_div/CryTmp[10][22] ), .CO(\u_div/CryTmp[10][23] ), 
        .S(\u_div/SumTmp[10][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_23  ( .A(\u_div/PartRem[11][23] ), .B(
        net31800), .CI(\u_div/CryTmp[10][23] ), .CO(\u_div/CryTmp[10][24] ), 
        .S(\u_div/SumTmp[10][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_19  ( .A(\u_div/PartRem[10][19] ), .B(
        net31910), .CI(\u_div/CryTmp[9][19] ), .CO(\u_div/CryTmp[9][20] ), .S(
        \u_div/SumTmp[9][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_1  ( .A(\u_div/PartRem[10][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[9][2] ), .S(
        \u_div/SumTmp[9][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_2  ( .A(\u_div/PartRem[10][2] ), .B(
        net32362), .CI(\u_div/CryTmp[9][2] ), .CO(\u_div/CryTmp[9][3] ), .S(
        \u_div/SumTmp[9][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_3  ( .A(\u_div/PartRem[10][3] ), .B(
        net32334), .CI(\u_div/CryTmp[9][3] ), .CO(\u_div/CryTmp[9][4] ), .S(
        \u_div/SumTmp[9][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_5  ( .A(\u_div/PartRem[10][5] ), .B(
        net32280), .CI(n768), .CO(\u_div/CryTmp[9][6] ), .S(
        \u_div/SumTmp[9][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_6  ( .A(\u_div/PartRem[10][6] ), .B(
        net32250), .CI(\u_div/CryTmp[9][6] ), .CO(\u_div/CryTmp[9][7] ), .S(
        \u_div/SumTmp[9][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_7  ( .A(\u_div/PartRem[10][7] ), .B(
        net32224), .CI(n316), .CO(\u_div/CryTmp[9][8] ), .S(
        \u_div/SumTmp[9][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_8  ( .A(\u_div/PartRem[10][8] ), .B(
        net32196), .CI(\u_div/CryTmp[9][8] ), .CO(\u_div/CryTmp[9][9] ), .S(
        \u_div/SumTmp[9][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_9  ( .A(\u_div/PartRem[10][9] ), .B(
        net32168), .CI(\u_div/CryTmp[9][9] ), .CO(\u_div/CryTmp[9][10] ), .S(
        \u_div/SumTmp[9][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_10  ( .A(\u_div/PartRem[10][10] ), .B(
        net32144), .CI(\u_div/CryTmp[9][10] ), .CO(\u_div/CryTmp[9][11] ), .S(
        \u_div/SumTmp[9][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_11  ( .A(\u_div/PartRem[10][11] ), .B(
        net32118), .CI(n302), .CO(\u_div/CryTmp[9][12] ), .S(
        \u_div/SumTmp[9][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_12  ( .A(\u_div/PartRem[10][12] ), .B(
        net32092), .CI(\u_div/CryTmp[9][12] ), .CO(\u_div/CryTmp[9][13] ), .S(
        \u_div/SumTmp[9][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_14  ( .A(\u_div/PartRem[10][14] ), .B(
        net32042), .CI(n187), .CO(\u_div/CryTmp[9][15] ), .S(
        \u_div/SumTmp[9][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_15  ( .A(\u_div/PartRem[10][15] ), .B(
        net32012), .CI(\u_div/CryTmp[9][15] ), .CO(\u_div/CryTmp[9][16] ), .S(
        \u_div/SumTmp[9][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_16  ( .A(\u_div/PartRem[10][16] ), .B(
        net31984), .CI(n139), .CO(\u_div/CryTmp[9][17] ), .S(
        \u_div/SumTmp[9][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_17  ( .A(\u_div/PartRem[10][17] ), .B(
        net31962), .CI(\u_div/CryTmp[9][17] ), .CO(\u_div/CryTmp[9][18] ), .S(
        \u_div/SumTmp[9][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_18  ( .A(\u_div/PartRem[10][18] ), .B(
        net31940), .CI(n113), .CO(\u_div/CryTmp[9][19] ), .S(
        \u_div/SumTmp[9][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_1  ( .A(\u_div/PartRem[9][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[8][2] ), .S(
        \u_div/SumTmp[8][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_2  ( .A(\u_div/PartRem[9][2] ), .B(
        net32362), .CI(\u_div/CryTmp[8][2] ), .CO(\u_div/CryTmp[8][3] ), .S(
        \u_div/SumTmp[8][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_3  ( .A(\u_div/CryTmp[8][3] ), .B(
        net32334), .CI(n244), .CO(\u_div/CryTmp[8][4] ), .S(
        \u_div/SumTmp[8][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_4  ( .A(\u_div/PartRem[9][4] ), .B(
        net32310), .CI(\u_div/CryTmp[8][4] ), .CO(\u_div/CryTmp[8][5] ), .S(
        \u_div/SumTmp[8][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_5  ( .A(\u_div/PartRem[9][5] ), .B(
        net32280), .CI(n119), .CO(\u_div/CryTmp[8][6] ), .S(
        \u_div/SumTmp[8][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_6  ( .A(\u_div/PartRem[9][6] ), .B(
        net32250), .CI(\u_div/CryTmp[8][6] ), .CO(\u_div/CryTmp[8][7] ), .S(
        \u_div/SumTmp[8][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_7  ( .A(\u_div/PartRem[9][7] ), .B(
        net32224), .CI(\u_div/CryTmp[8][7] ), .CO(\u_div/CryTmp[8][8] ), .S(
        \u_div/SumTmp[8][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_8  ( .A(\u_div/PartRem[9][8] ), .B(
        net32196), .CI(n2), .CO(\u_div/CryTmp[8][9] ), .S(\u_div/SumTmp[8][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_9  ( .A(\u_div/PartRem[9][9] ), .B(
        net32168), .CI(\u_div/CryTmp[8][9] ), .CO(\u_div/CryTmp[8][10] ), .S(
        \u_div/SumTmp[8][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_10  ( .A(\u_div/PartRem[9][10] ), .B(
        net32144), .CI(n772), .CO(\u_div/CryTmp[8][11] ), .S(
        \u_div/SumTmp[8][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_11  ( .A(\u_div/PartRem[9][11] ), .B(
        net32118), .CI(n774), .CO(\u_div/CryTmp[8][12] ), .S(
        \u_div/SumTmp[8][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_12  ( .A(\u_div/PartRem[9][12] ), .B(
        \u_div/CryTmp[8][12] ), .CI(net32092), .CO(\u_div/CryTmp[8][13] ), .S(
        \u_div/SumTmp[8][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_14  ( .A(\u_div/PartRem[9][14] ), .B(
        net32042), .CI(n770), .CO(\u_div/CryTmp[8][15] ), .S(
        \u_div/SumTmp[8][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_15  ( .A(\u_div/PartRem[9][15] ), .B(
        net32012), .CI(\u_div/CryTmp[8][15] ), .CO(\u_div/CryTmp[8][16] ), .S(
        \u_div/SumTmp[8][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_16  ( .A(\u_div/PartRem[9][16] ), .B(
        net31984), .CI(\u_div/CryTmp[8][16] ), .CO(\u_div/CryTmp[8][17] ), .S(
        \u_div/SumTmp[8][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_17  ( .A(\u_div/PartRem[9][17] ), .B(
        net31962), .CI(\u_div/CryTmp[8][17] ), .CO(\u_div/CryTmp[8][18] ), .S(
        \u_div/SumTmp[8][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_18  ( .A(\u_div/PartRem[9][18] ), .B(
        net31940), .CI(\u_div/CryTmp[8][18] ), .CO(\u_div/CryTmp[8][19] ), .S(
        \u_div/SumTmp[8][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_19  ( .A(\u_div/PartRem[9][19] ), .B(
        net31910), .CI(\u_div/CryTmp[8][19] ), .CO(\u_div/CryTmp[8][20] ), .S(
        \u_div/SumTmp[8][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_7_20  ( .A(\u_div/PartRem[8][20] ), .B(
        net31882), .CI(\u_div/CryTmp[7][20] ), .CO(\u_div/CryTmp[7][21] ), .S(
        \u_div/SumTmp[7][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_20  ( .A(\u_div/PartRem[15][20] ), .B(
        net31884), .CI(\u_div/CryTmp[14][20] ), .CO(\u_div/CryTmp[14][21] ), 
        .S(\u_div/SumTmp[14][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_1  ( .A(n758), .B(net32384), .CI(
        \u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[14][2] ), .S(
        \u_div/SumTmp[14][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_2  ( .A(\u_div/PartRem[15][2] ), .B(
        net32364), .CI(\u_div/CryTmp[14][2] ), .CO(\u_div/CryTmp[14][3] ), .S(
        \u_div/SumTmp[14][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_3  ( .A(\u_div/PartRem[15][3] ), .B(
        net32336), .CI(\u_div/CryTmp[14][3] ), .CO(\u_div/CryTmp[14][4] ), .S(
        \u_div/SumTmp[14][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_4  ( .A(\u_div/PartRem[15][4] ), .B(
        net32312), .CI(\u_div/CryTmp[14][4] ), .CO(\u_div/CryTmp[14][5] ), .S(
        \u_div/SumTmp[14][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_5  ( .A(\u_div/PartRem[15][5] ), .B(
        net32282), .CI(\u_div/CryTmp[14][5] ), .CO(\u_div/CryTmp[14][6] ), .S(
        \u_div/SumTmp[14][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_6  ( .A(\u_div/PartRem[15][6] ), .B(
        net32252), .CI(\u_div/CryTmp[14][6] ), .CO(\u_div/CryTmp[14][7] ), .S(
        \u_div/SumTmp[14][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_7  ( .A(\u_div/PartRem[15][7] ), .B(
        net32224), .CI(\u_div/CryTmp[14][7] ), .CO(\u_div/CryTmp[14][8] ), .S(
        \u_div/SumTmp[14][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_8  ( .A(\u_div/PartRem[15][8] ), .B(
        net32198), .CI(\u_div/CryTmp[14][8] ), .CO(\u_div/CryTmp[14][9] ), .S(
        \u_div/SumTmp[14][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_9  ( .A(\u_div/PartRem[15][9] ), .B(
        net32166), .CI(\u_div/CryTmp[14][9] ), .CO(\u_div/CryTmp[14][10] ), 
        .S(\u_div/SumTmp[14][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_10  ( .A(\u_div/PartRem[15][10] ), .B(
        net32142), .CI(\u_div/CryTmp[14][10] ), .CO(\u_div/CryTmp[14][11] ), 
        .S(\u_div/SumTmp[14][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_11  ( .A(\u_div/PartRem[15][11] ), .B(
        net32116), .CI(\u_div/CryTmp[14][11] ), .CO(\u_div/CryTmp[14][12] ), 
        .S(\u_div/SumTmp[14][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_13  ( .A(\u_div/PartRem[15][13] ), .B(
        net32066), .CI(\u_div/CryTmp[14][13] ), .CO(\u_div/CryTmp[14][14] ), 
        .S(\u_div/SumTmp[14][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_14  ( .A(\u_div/PartRem[15][14] ), .B(
        net32044), .CI(\u_div/CryTmp[14][14] ), .CO(\u_div/CryTmp[14][15] ), 
        .S(\u_div/SumTmp[14][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_16  ( .A(\u_div/PartRem[15][16] ), .B(
        net31984), .CI(n747), .CO(\u_div/CryTmp[14][17] ), .S(
        \u_div/SumTmp[14][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_17  ( .A(\u_div/PartRem[15][17] ), .B(
        net31962), .CI(\u_div/CryTmp[14][17] ), .CO(\u_div/CryTmp[14][18] ), 
        .S(\u_div/SumTmp[14][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_18  ( .A(\u_div/PartRem[15][18] ), .B(
        net31940), .CI(n117), .CO(\u_div/CryTmp[14][19] ), .S(
        \u_div/SumTmp[14][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_19  ( .A(\u_div/PartRem[15][19] ), .B(
        net31912), .CI(\u_div/CryTmp[14][19] ), .CO(\u_div/CryTmp[14][20] ), 
        .S(\u_div/SumTmp[14][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_1  ( .A(\u_div/PartRem[14][1] ), .B(
        net32384), .CI(\u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[13][2] ), .S(
        \u_div/SumTmp[13][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_2  ( .A(\u_div/PartRem[14][2] ), .B(
        net32364), .CI(\u_div/CryTmp[13][2] ), .CO(\u_div/CryTmp[13][3] ), .S(
        \u_div/SumTmp[13][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_3  ( .A(\u_div/PartRem[14][3] ), .B(
        net32336), .CI(\u_div/CryTmp[13][3] ), .CO(\u_div/CryTmp[13][4] ), .S(
        \u_div/SumTmp[13][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_4  ( .A(\u_div/PartRem[14][4] ), .B(
        net32312), .CI(\u_div/CryTmp[13][4] ), .CO(\u_div/CryTmp[13][5] ), .S(
        \u_div/SumTmp[13][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_5  ( .A(\u_div/PartRem[14][5] ), .B(
        net32282), .CI(\u_div/CryTmp[13][5] ), .CO(\u_div/CryTmp[13][6] ), .S(
        \u_div/SumTmp[13][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_6  ( .A(\u_div/PartRem[14][6] ), .B(
        net32252), .CI(\u_div/CryTmp[13][6] ), .CO(\u_div/CryTmp[13][7] ), .S(
        \u_div/SumTmp[13][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_7  ( .A(n189), .B(net32224), .CI(
        \u_div/CryTmp[13][7] ), .CO(\u_div/CryTmp[13][8] ), .S(
        \u_div/SumTmp[13][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_8  ( .A(\u_div/PartRem[14][8] ), .B(
        net32198), .CI(\u_div/CryTmp[13][8] ), .CO(\u_div/CryTmp[13][9] ), .S(
        \u_div/SumTmp[13][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_9  ( .A(\u_div/PartRem[14][9] ), .B(
        net32168), .CI(\u_div/CryTmp[13][9] ), .CO(\u_div/CryTmp[13][10] ), 
        .S(\u_div/SumTmp[13][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_10  ( .A(n31), .B(net32142), .CI(n83), 
        .CO(\u_div/CryTmp[13][11] ), .S(\u_div/SumTmp[13][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_11  ( .A(\u_div/PartRem[14][11] ), .B(
        net32116), .CI(\u_div/CryTmp[13][11] ), .CO(\u_div/CryTmp[13][12] ), 
        .S(\u_div/SumTmp[13][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_12  ( .A(\u_div/PartRem[14][12] ), .B(
        net32090), .CI(\u_div/CryTmp[13][12] ), .CO(\u_div/CryTmp[13][13] ), 
        .S(\u_div/SumTmp[13][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_13  ( .A(\u_div/PartRem[14][13] ), .B(
        net32066), .CI(\u_div/CryTmp[13][13] ), .CO(\u_div/CryTmp[13][14] ), 
        .S(\u_div/SumTmp[13][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_14  ( .A(\u_div/PartRem[14][14] ), .B(
        net32044), .CI(\u_div/CryTmp[13][14] ), .CO(\u_div/CryTmp[13][15] ), 
        .S(\u_div/SumTmp[13][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_15  ( .A(\u_div/PartRem[14][15] ), .B(
        net32014), .CI(\u_div/CryTmp[13][15] ), .CO(\u_div/CryTmp[13][16] ), 
        .S(\u_div/SumTmp[13][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_16  ( .A(\u_div/PartRem[14][16] ), .B(
        net31984), .CI(\u_div/CryTmp[13][16] ), .CO(\u_div/CryTmp[13][17] ), 
        .S(\u_div/SumTmp[13][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_18  ( .A(\u_div/PartRem[14][18] ), .B(
        net31940), .CI(n739), .CO(\u_div/CryTmp[13][19] ), .S(
        \u_div/SumTmp[13][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_19  ( .A(\u_div/PartRem[14][19] ), .B(
        net31912), .CI(\u_div/CryTmp[13][19] ), .CO(\u_div/CryTmp[13][20] ), 
        .S(\u_div/SumTmp[13][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_20  ( .A(\u_div/PartRem[14][20] ), .B(
        net31884), .CI(\u_div/CryTmp[13][20] ), .CO(\u_div/CryTmp[13][21] ), 
        .S(\u_div/SumTmp[13][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_12  ( .A(\u_div/PartRem[12][12] ), .B(
        net32090), .CI(n754), .CO(\u_div/CryTmp[11][13] ), .S(
        \u_div/SumTmp[11][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_13  ( .A(n99), .B(net32066), .CI(
        \u_div/CryTmp[11][13] ), .CO(\u_div/CryTmp[11][14] ), .S(
        \u_div/SumTmp[11][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_14  ( .A(\u_div/PartRem[12][14] ), .B(
        net32042), .CI(\u_div/CryTmp[11][14] ), .CO(\u_div/CryTmp[11][15] ), 
        .S(\u_div/SumTmp[11][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_15  ( .A(\u_div/PartRem[12][15] ), .B(
        net32012), .CI(\u_div/CryTmp[11][15] ), .CO(\u_div/CryTmp[11][16] ), 
        .S(\u_div/SumTmp[11][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_16  ( .A(\u_div/PartRem[12][16] ), .B(
        net31984), .CI(\u_div/CryTmp[11][16] ), .CO(\u_div/CryTmp[11][17] ), 
        .S(\u_div/SumTmp[11][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_17  ( .A(\u_div/PartRem[12][17] ), .B(
        net31962), .CI(n36), .CO(\u_div/CryTmp[11][18] ), .S(
        \u_div/SumTmp[11][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_19  ( .A(net31910), .B(n749), .CI(
        \u_div/PartRem[12][19] ), .CO(\u_div/CryTmp[11][20] ), .S(
        \u_div/SumTmp[11][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_20  ( .A(\u_div/PartRem[12][20] ), .B(
        net31882), .CI(n312), .CO(\u_div/CryTmp[11][21] ), .S(
        \u_div/SumTmp[11][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_21  ( .A(\u_div/PartRem[12][21] ), .B(
        net31854), .CI(\u_div/CryTmp[11][21] ), .CO(\u_div/CryTmp[11][22] ), 
        .S(\u_div/SumTmp[11][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_22  ( .A(\u_div/PartRem[12][22] ), .B(
        net31826), .CI(\u_div/CryTmp[11][22] ), .CO(\u_div/CryTmp[11][23] ), 
        .S(\u_div/SumTmp[11][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_23  ( .A(\u_div/PartRem[12][23] ), .B(
        net31800), .CI(n105), .CO(\u_div/CryTmp[11][24] ), .S(
        \u_div/SumTmp[11][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_1  ( .A(\u_div/PartRem[13][1] ), .B(
        net32384), .CI(\u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[12][2] ), .S(
        \u_div/SumTmp[12][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_2  ( .A(\u_div/PartRem[13][2] ), .B(
        net32364), .CI(\u_div/CryTmp[12][2] ), .CO(\u_div/CryTmp[12][3] ), .S(
        \u_div/SumTmp[12][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_3  ( .A(\u_div/PartRem[13][3] ), .B(
        net32336), .CI(\u_div/CryTmp[12][3] ), .CO(\u_div/CryTmp[12][4] ), .S(
        \u_div/SumTmp[12][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_4  ( .A(\u_div/PartRem[13][4] ), .B(
        net32312), .CI(\u_div/CryTmp[12][4] ), .CO(\u_div/CryTmp[12][5] ), .S(
        \u_div/SumTmp[12][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_5  ( .A(\u_div/PartRem[13][5] ), .B(
        net32282), .CI(\u_div/CryTmp[12][5] ), .CO(\u_div/CryTmp[12][6] ), .S(
        \u_div/SumTmp[12][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_6  ( .A(\u_div/PartRem[13][6] ), .B(
        net32252), .CI(\u_div/CryTmp[12][6] ), .CO(\u_div/CryTmp[12][7] ), .S(
        \u_div/SumTmp[12][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_7  ( .A(\u_div/PartRem[13][7] ), .B(
        net32224), .CI(\u_div/CryTmp[12][7] ), .CO(\u_div/CryTmp[12][8] ), .S(
        \u_div/SumTmp[12][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_8  ( .A(\u_div/PartRem[13][8] ), .B(
        net32198), .CI(\u_div/CryTmp[12][8] ), .CO(\u_div/CryTmp[12][9] ), .S(
        \u_div/SumTmp[12][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_9  ( .A(\u_div/PartRem[13][9] ), .B(
        net32168), .CI(\u_div/CryTmp[12][9] ), .CO(\u_div/CryTmp[12][10] ), 
        .S(\u_div/SumTmp[12][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_10  ( .A(n81), .B(net32144), .CI(
        \u_div/CryTmp[12][10] ), .CO(\u_div/CryTmp[12][11] ), .S(
        \u_div/SumTmp[12][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_11  ( .A(\u_div/PartRem[13][11] ), .B(
        net32116), .CI(\u_div/CryTmp[12][11] ), .CO(\u_div/CryTmp[12][12] ), 
        .S(\u_div/SumTmp[12][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_12  ( .A(\u_div/PartRem[13][12] ), .B(
        net32090), .CI(\u_div/CryTmp[12][12] ), .CO(\u_div/CryTmp[12][13] ), 
        .S(\u_div/SumTmp[12][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_13  ( .A(\u_div/PartRem[13][13] ), .B(
        net32066), .CI(\u_div/CryTmp[12][13] ), .CO(\u_div/CryTmp[12][14] ), 
        .S(\u_div/SumTmp[12][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_14  ( .A(\u_div/PartRem[13][14] ), .B(
        net32044), .CI(\u_div/CryTmp[12][14] ), .CO(\u_div/CryTmp[12][15] ), 
        .S(\u_div/SumTmp[12][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_16  ( .A(net31984), .B(
        \u_div/PartRem[13][16] ), .CI(\u_div/CryTmp[12][16] ), .CO(
        \u_div/CryTmp[12][17] ), .S(\u_div/SumTmp[12][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_17  ( .A(net31962), .B(
        \u_div/PartRem[13][17] ), .CI(\u_div/CryTmp[12][17] ), .CO(
        \u_div/CryTmp[12][18] ), .S(\u_div/SumTmp[12][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_19  ( .A(\u_div/PartRem[13][19] ), .B(
        net31912), .CI(n760), .CO(\u_div/CryTmp[12][20] ), .S(
        \u_div/SumTmp[12][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_22  ( .A(\u_div/PartRem[13][22] ), .B(
        net31828), .CI(n741), .CO(\u_div/CryTmp[12][23] ), .S(
        \u_div/SumTmp[12][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_23  ( .A(\u_div/PartRem[13][23] ), .B(
        net31802), .CI(n743), .CO(\u_div/CryTmp[12][24] ), .S(
        \u_div/SumTmp[12][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_1  ( .A(\u_div/PartRem[12][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[11][2] ), .S(
        \u_div/SumTmp[11][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_2  ( .A(\u_div/PartRem[12][2] ), .B(
        net32362), .CI(\u_div/CryTmp[11][2] ), .CO(\u_div/CryTmp[11][3] ), .S(
        \u_div/SumTmp[11][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_3  ( .A(\u_div/PartRem[12][3] ), .B(
        net32334), .CI(\u_div/CryTmp[11][3] ), .CO(\u_div/CryTmp[11][4] ), .S(
        \u_div/SumTmp[11][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_4  ( .A(\u_div/PartRem[12][4] ), .B(
        net32310), .CI(\u_div/CryTmp[11][4] ), .CO(\u_div/CryTmp[11][5] ), .S(
        \u_div/SumTmp[11][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_5  ( .A(\u_div/PartRem[12][5] ), .B(
        net32280), .CI(\u_div/CryTmp[11][5] ), .CO(\u_div/CryTmp[11][6] ), .S(
        \u_div/SumTmp[11][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_6  ( .A(\u_div/PartRem[12][6] ), .B(
        net32250), .CI(\u_div/CryTmp[11][6] ), .CO(\u_div/CryTmp[11][7] ), .S(
        \u_div/SumTmp[11][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_7  ( .A(\u_div/PartRem[12][7] ), .B(
        net32224), .CI(\u_div/CryTmp[11][7] ), .CO(\u_div/CryTmp[11][8] ), .S(
        \u_div/SumTmp[11][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_8  ( .A(\u_div/PartRem[12][8] ), .B(
        net32196), .CI(\u_div/CryTmp[11][8] ), .CO(\u_div/CryTmp[11][9] ), .S(
        \u_div/SumTmp[11][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_10  ( .A(\u_div/PartRem[12][10] ), .B(
        net32144), .CI(n109), .CO(\u_div/CryTmp[11][11] ), .S(
        \u_div/SumTmp[11][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_11  ( .A(net45940), .B(net32118), .CI(
        \u_div/CryTmp[11][11] ), .CO(\u_div/CryTmp[11][12] ), .S(
        \u_div/SumTmp[11][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_1  ( .A(\u_div/PartRem[11][1] ), .B(
        net32382), .CI(\u_div/CryTmp[11][1] ), .CO(\u_div/CryTmp[10][2] ), .S(
        \u_div/SumTmp[10][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_2  ( .A(\u_div/PartRem[11][2] ), .B(
        net32362), .CI(\u_div/CryTmp[10][2] ), .CO(\u_div/CryTmp[10][3] ), .S(
        \u_div/SumTmp[10][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_3  ( .A(\u_div/PartRem[11][3] ), .B(
        net32334), .CI(\u_div/CryTmp[10][3] ), .CO(\u_div/CryTmp[10][4] ), .S(
        \u_div/SumTmp[10][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_4  ( .A(\u_div/PartRem[11][4] ), .B(
        net32310), .CI(\u_div/CryTmp[10][4] ), .CO(\u_div/CryTmp[10][5] ), .S(
        \u_div/SumTmp[10][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_5  ( .A(\u_div/PartRem[11][5] ), .B(
        net32280), .CI(\u_div/CryTmp[10][5] ), .CO(\u_div/CryTmp[10][6] ), .S(
        \u_div/SumTmp[10][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_6  ( .A(\u_div/PartRem[11][6] ), .B(
        net32250), .CI(\u_div/CryTmp[10][6] ), .CO(\u_div/CryTmp[10][7] ), .S(
        \u_div/SumTmp[10][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_7  ( .A(\u_div/PartRem[11][7] ), .B(
        net32224), .CI(\u_div/CryTmp[10][7] ), .CO(\u_div/CryTmp[10][8] ), .S(
        \u_div/SumTmp[10][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_8  ( .A(\u_div/PartRem[11][8] ), .B(
        net32196), .CI(\u_div/CryTmp[10][8] ), .CO(\u_div/CryTmp[10][9] ), .S(
        \u_div/SumTmp[10][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_9  ( .A(\u_div/PartRem[11][9] ), .B(
        net32168), .CI(\u_div/CryTmp[10][9] ), .CO(\u_div/CryTmp[10][10] ), 
        .S(\u_div/SumTmp[10][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_10  ( .A(\u_div/PartRem[11][10] ), .B(
        net32144), .CI(\u_div/CryTmp[10][10] ), .CO(\u_div/CryTmp[10][11] ), 
        .S(\u_div/SumTmp[10][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_11  ( .A(n751), .B(net32118), .CI(n745), 
        .CO(\u_div/CryTmp[10][12] ), .S(\u_div/SumTmp[10][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_12  ( .A(net46752), .B(net32092), .CI(
        n756), .CO(\u_div/CryTmp[10][13] ), .S(\u_div/SumTmp[10][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_13  ( .A(\u_div/PartRem[11][13] ), .B(
        net32066), .CI(\u_div/CryTmp[10][13] ), .CO(\u_div/CryTmp[10][14] ), 
        .S(\u_div/SumTmp[10][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_14  ( .A(\u_div/PartRem[11][14] ), .B(
        net32042), .CI(\u_div/CryTmp[10][14] ), .CO(\u_div/CryTmp[10][15] ), 
        .S(\u_div/SumTmp[10][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_15  ( .A(\u_div/PartRem[11][15] ), .B(
        net32012), .CI(n306), .CO(\u_div/CryTmp[10][16] ), .S(
        \u_div/SumTmp[10][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_2  ( .A(\u_div/PartRem[17][2] ), .B(
        net32364), .CI(\u_div/CryTmp[16][2] ), .CO(\u_div/CryTmp[16][3] ), .S(
        \u_div/SumTmp[16][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_3  ( .A(\u_div/PartRem[17][3] ), .B(
        net32336), .CI(n290), .CO(\u_div/CryTmp[16][4] ), .S(
        \u_div/SumTmp[16][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_5  ( .A(\u_div/PartRem[17][5] ), .B(
        net32282), .CI(n288), .CO(\u_div/CryTmp[16][6] ), .S(
        \u_div/SumTmp[16][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_6  ( .A(\u_div/PartRem[17][6] ), .B(
        net32252), .CI(\u_div/CryTmp[16][6] ), .CO(\u_div/CryTmp[16][7] ), .S(
        \u_div/SumTmp[16][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_7  ( .A(\u_div/PartRem[17][7] ), .B(
        net32222), .CI(n155), .CO(\u_div/CryTmp[16][8] ), .S(
        \u_div/SumTmp[16][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_8  ( .A(\u_div/PartRem[17][8] ), .B(
        net32198), .CI(\u_div/CryTmp[16][8] ), .CO(\u_div/CryTmp[16][9] ), .S(
        \u_div/SumTmp[16][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_9  ( .A(\u_div/PartRem[17][9] ), .B(
        net32166), .CI(\u_div/CryTmp[16][9] ), .CO(\u_div/CryTmp[16][10] ), 
        .S(\u_div/SumTmp[16][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_10  ( .A(\u_div/PartRem[17][10] ), .B(
        net32142), .CI(\u_div/CryTmp[16][10] ), .CO(\u_div/CryTmp[16][11] ), 
        .S(\u_div/SumTmp[16][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_11  ( .A(\u_div/PartRem[17][11] ), .B(
        net32116), .CI(\u_div/CryTmp[16][11] ), .CO(\u_div/CryTmp[16][12] ), 
        .S(\u_div/SumTmp[16][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_12  ( .A(\u_div/PartRem[17][12] ), .B(
        net32090), .CI(\u_div/CryTmp[16][12] ), .CO(\u_div/CryTmp[16][13] ), 
        .S(\u_div/SumTmp[16][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_13  ( .A(\u_div/PartRem[17][13] ), .B(
        net32066), .CI(n44), .CO(\u_div/CryTmp[16][14] ), .S(
        \u_div/SumTmp[16][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_14  ( .A(\u_div/PartRem[17][14] ), .B(
        net32044), .CI(\u_div/CryTmp[16][14] ), .CO(\u_div/CryTmp[16][15] ), 
        .S(\u_div/SumTmp[16][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_15  ( .A(\u_div/PartRem[17][15] ), .B(
        net32014), .CI(n677), .CO(\u_div/CryTmp[16][16] ), .S(
        \u_div/SumTmp[16][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_16  ( .A(\u_div/PartRem[17][16] ), .B(
        net31984), .CI(\u_div/CryTmp[16][16] ), .CO(\u_div/CryTmp[16][17] ), 
        .S(\u_div/SumTmp[16][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_17  ( .A(\u_div/PartRem[17][17] ), .B(
        net31962), .CI(\u_div/CryTmp[16][17] ), .CO(\u_div/CryTmp[16][18] ), 
        .S(\u_div/SumTmp[16][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_18  ( .A(net31938), .B(
        \u_div/PartRem[17][18] ), .CI(n131), .CO(\u_div/CryTmp[16][19] ), .S(
        \u_div/SumTmp[16][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_19  ( .A(\u_div/PartRem[17][19] ), .B(
        net31912), .CI(\u_div/CryTmp[16][19] ), .CO(\u_div/CryTmp[16][20] ), 
        .S(\u_div/SumTmp[16][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_20  ( .A(\u_div/PartRem[17][20] ), .B(
        net31884), .CI(\u_div/CryTmp[16][20] ), .CO(\u_div/CryTmp[16][21] ), 
        .S(\u_div/SumTmp[16][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_21  ( .A(net52402), .B(net31856), .CI(
        n680), .CO(\u_div/CryTmp[16][22] ), .S(\u_div/SumTmp[16][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_22  ( .A(\u_div/PartRem[17][22] ), .B(
        net31828), .CI(\u_div/CryTmp[16][22] ), .CO(\u_div/CryTmp[16][23] ), 
        .S(\u_div/SumTmp[16][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_23  ( .A(\u_div/PartRem[17][23] ), .B(
        net31802), .CI(n97), .CO(\u_div/CryTmp[16][24] ), .S(
        \u_div/SumTmp[16][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_12  ( .A(\u_div/PartRem[16][12] ), .B(
        net32090), .CI(n298), .CO(\u_div/CryTmp[15][13] ), .S(
        \u_div/SumTmp[15][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_13  ( .A(\u_div/PartRem[16][13] ), .B(
        net32066), .CI(\u_div/CryTmp[15][13] ), .CO(\u_div/CryTmp[15][14] ), 
        .S(\u_div/SumTmp[15][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_14  ( .A(\u_div/PartRem[16][14] ), .B(
        net32044), .CI(\u_div/CryTmp[15][14] ), .CO(\u_div/CryTmp[15][15] ), 
        .S(\u_div/SumTmp[15][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_15  ( .A(\u_div/PartRem[16][15] ), .B(
        net32014), .CI(\u_div/CryTmp[15][15] ), .CO(\u_div/CryTmp[15][16] ), 
        .S(\u_div/SumTmp[15][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_16  ( .A(n101), .B(net31984), .CI(
        \u_div/PartRem[16][16] ), .CO(\u_div/CryTmp[15][17] ), .S(
        \u_div/SumTmp[15][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_17  ( .A(\u_div/PartRem[16][17] ), .B(
        net31962), .CI(\u_div/CryTmp[15][17] ), .CO(\u_div/CryTmp[15][18] ), 
        .S(\u_div/SumTmp[15][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_18  ( .A(\u_div/PartRem[16][18] ), .B(
        net31940), .CI(\u_div/CryTmp[15][18] ), .CO(\u_div/CryTmp[15][19] ), 
        .S(\u_div/SumTmp[15][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_20  ( .A(\u_div/PartRem[16][20] ), .B(
        n320), .CI(net31884), .CO(\u_div/CryTmp[15][21] ), .S(
        \u_div/SumTmp[15][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_21  ( .A(\u_div/PartRem[16][21] ), .B(
        net31856), .CI(n318), .CO(\u_div/CryTmp[15][22] ), .S(
        \u_div/SumTmp[15][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_22  ( .A(\u_div/PartRem[16][22] ), .B(
        net31828), .CI(\u_div/CryTmp[15][22] ), .CO(\u_div/CryTmp[15][23] ), 
        .S(\u_div/SumTmp[15][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_23  ( .A(\u_div/PartRem[16][23] ), .B(
        net31802), .CI(\u_div/CryTmp[15][23] ), .CO(\u_div/CryTmp[15][24] ), 
        .S(\u_div/SumTmp[15][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_1  ( .A(\u_div/PartRem[16][1] ), .B(
        net32384), .CI(\u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[15][2] ), .S(
        \u_div/SumTmp[15][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_2  ( .A(\u_div/PartRem[16][2] ), .B(
        net32364), .CI(\u_div/CryTmp[15][2] ), .CO(\u_div/CryTmp[15][3] ), .S(
        \u_div/SumTmp[15][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_3  ( .A(\u_div/PartRem[16][3] ), .B(
        net32336), .CI(n24), .CO(\u_div/CryTmp[15][4] ), .S(
        \u_div/SumTmp[15][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_4  ( .A(\u_div/PartRem[16][4] ), .B(
        net32312), .CI(\u_div/CryTmp[15][4] ), .CO(\u_div/CryTmp[15][5] ), .S(
        \u_div/SumTmp[15][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_5  ( .A(\u_div/CryTmp[15][5] ), .B(
        net32282), .CI(\u_div/PartRem[16][5] ), .CO(\u_div/CryTmp[15][6] ), 
        .S(\u_div/SumTmp[15][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_6  ( .A(\u_div/PartRem[16][6] ), .B(
        net32252), .CI(\u_div/CryTmp[15][6] ), .CO(\u_div/CryTmp[15][7] ), .S(
        \u_div/SumTmp[15][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_7  ( .A(\u_div/PartRem[16][7] ), .B(
        net32224), .CI(\u_div/CryTmp[15][7] ), .CO(\u_div/CryTmp[15][8] ), .S(
        \u_div/SumTmp[15][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_8  ( .A(\u_div/PartRem[16][8] ), .B(
        net32198), .CI(\u_div/CryTmp[15][8] ), .CO(\u_div/CryTmp[15][9] ), .S(
        \u_div/SumTmp[15][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_9  ( .A(\u_div/PartRem[16][9] ), .B(
        net32166), .CI(\u_div/CryTmp[15][9] ), .CO(\u_div/CryTmp[15][10] ), 
        .S(\u_div/SumTmp[15][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_10  ( .A(\u_div/PartRem[16][10] ), .B(
        net32142), .CI(\u_div/CryTmp[15][10] ), .CO(\u_div/CryTmp[15][11] ), 
        .S(\u_div/SumTmp[15][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_14_12  ( .A(\u_div/PartRem[15][12] ), .B(
        net32090), .CI(net42406), .CO(\u_div/CryTmp[14][13] ), .S(
        \u_div/SumTmp[14][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_18  ( .A(\u_div/PartRem[21][18] ), .B(
        net31938), .CI(n63), .CO(\u_div/CryTmp[20][19] ), .S(
        \u_div/SumTmp[20][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_19  ( .A(\u_div/PartRem[21][19] ), .B(
        net31912), .CI(\u_div/CryTmp[20][19] ), .CO(\u_div/CryTmp[20][20] ), 
        .S(\u_div/SumTmp[20][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_20  ( .A(\u_div/PartRem[21][20] ), .B(
        net31884), .CI(\u_div/CryTmp[20][20] ), .CO(\u_div/CryTmp[20][21] ), 
        .S(\u_div/SumTmp[20][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_21  ( .A(\u_div/PartRem[21][21] ), .B(
        net31856), .CI(\u_div/CryTmp[20][21] ), .CO(\u_div/CryTmp[20][22] ), 
        .S(\u_div/SumTmp[20][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_22  ( .A(\u_div/PartRem[21][22] ), .B(
        net31828), .CI(n644), .CO(\u_div/CryTmp[20][23] ), .S(
        \u_div/SumTmp[20][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_23  ( .A(\u_div/PartRem[21][23] ), .B(
        net31802), .CI(\u_div/CryTmp[20][23] ), .CO(\u_div/CryTmp[20][24] ), 
        .S(\u_div/SumTmp[20][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_19  ( .A(\u_div/PartRem[20][19] ), .B(
        net31912), .CI(\u_div/CryTmp[19][19] ), .CO(\u_div/CryTmp[19][20] ), 
        .S(\u_div/SumTmp[19][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_20  ( .A(\u_div/PartRem[20][20] ), .B(
        net31884), .CI(\u_div/CryTmp[19][20] ), .CO(\u_div/CryTmp[19][21] ), 
        .S(\u_div/SumTmp[19][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_21  ( .A(\u_div/PartRem[20][21] ), .B(
        net31856), .CI(\u_div/CryTmp[19][21] ), .CO(\u_div/CryTmp[19][22] ), 
        .S(\u_div/SumTmp[19][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_22  ( .A(\u_div/PartRem[20][22] ), .B(
        net31828), .CI(\u_div/CryTmp[19][22] ), .CO(\u_div/CryTmp[19][23] ), 
        .S(\u_div/SumTmp[19][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_23  ( .A(\u_div/PartRem[20][23] ), .B(
        net31802), .CI(\u_div/CryTmp[19][23] ), .CO(\u_div/CryTmp[19][24] ), 
        .S(\u_div/SumTmp[19][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_1  ( .A(\u_div/PartRem[18][1] ), .B(
        net32384), .CI(\u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[17][2] ), .S(
        \u_div/SumTmp[17][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_2  ( .A(\u_div/PartRem[18][2] ), .B(
        net32364), .CI(n256), .CO(\u_div/CryTmp[17][3] ), .S(
        \u_div/SumTmp[17][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_3  ( .A(\u_div/PartRem[18][3] ), .B(
        net32336), .CI(\u_div/CryTmp[17][3] ), .CO(\u_div/CryTmp[17][4] ), .S(
        \u_div/SumTmp[17][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_4  ( .A(\u_div/PartRem[18][4] ), .B(
        net32312), .CI(\u_div/CryTmp[17][4] ), .CO(\u_div/CryTmp[17][5] ), .S(
        \u_div/SumTmp[17][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_5  ( .A(\u_div/PartRem[18][5] ), .B(
        net32282), .CI(\u_div/CryTmp[17][5] ), .CO(\u_div/CryTmp[17][6] ), .S(
        \u_div/SumTmp[17][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_8  ( .A(\u_div/PartRem[18][8] ), .B(
        net32198), .CI(n640), .CO(\u_div/CryTmp[17][9] ), .S(
        \u_div/SumTmp[17][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_9  ( .A(\u_div/PartRem[18][9] ), .B(
        net32166), .CI(\u_div/CryTmp[17][9] ), .CO(\u_div/CryTmp[17][10] ), 
        .S(\u_div/SumTmp[17][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_10  ( .A(\u_div/PartRem[18][10] ), .B(
        net32142), .CI(\u_div/CryTmp[17][10] ), .CO(\u_div/CryTmp[17][11] ), 
        .S(\u_div/SumTmp[17][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_11  ( .A(\u_div/PartRem[18][11] ), .B(
        net32116), .CI(\u_div/CryTmp[17][11] ), .CO(\u_div/CryTmp[17][12] ), 
        .S(\u_div/SumTmp[17][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_12  ( .A(\u_div/PartRem[18][12] ), .B(
        \u_div/CryTmp[17][12] ), .CI(net32090), .CO(\u_div/CryTmp[17][13] ), 
        .S(\u_div/SumTmp[17][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_13  ( .A(\u_div/PartRem[18][13] ), .B(
        net32066), .CI(\u_div/CryTmp[17][13] ), .CO(\u_div/CryTmp[17][14] ), 
        .S(\u_div/SumTmp[17][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_14  ( .A(\u_div/PartRem[18][14] ), .B(
        net32044), .CI(n630), .CO(\u_div/CryTmp[17][15] ), .S(
        \u_div/SumTmp[17][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_15  ( .A(\u_div/PartRem[18][15] ), .B(
        net32014), .CI(\u_div/CryTmp[17][15] ), .CO(\u_div/CryTmp[17][16] ), 
        .S(\u_div/SumTmp[17][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_16  ( .A(\u_div/PartRem[18][16] ), .B(
        net31984), .CI(\u_div/CryTmp[17][16] ), .CO(\u_div/CryTmp[17][17] ), 
        .S(\u_div/SumTmp[17][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_17  ( .A(\u_div/PartRem[18][17] ), .B(
        net31962), .CI(\u_div/CryTmp[17][17] ), .CO(\u_div/CryTmp[17][18] ), 
        .S(\u_div/SumTmp[17][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_19  ( .A(\u_div/PartRem[18][19] ), .B(
        net31912), .CI(n632), .CO(\u_div/CryTmp[17][20] ), .S(
        \u_div/SumTmp[17][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_20  ( .A(n642), .B(net31884), .CI(
        \u_div/PartRem[18][20] ), .CO(\u_div/CryTmp[17][21] ), .S(
        \u_div/SumTmp[17][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_22  ( .A(n296), .B(net31828), .CI(
        \u_div/PartRem[18][22] ), .CO(\u_div/CryTmp[17][23] ), .S(
        \u_div/SumTmp[17][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_23  ( .A(n638), .B(net31802), .CI(
        \u_div/CryTmp[17][23] ), .CO(\u_div/CryTmp[17][24] ), .S(
        \u_div/SumTmp[17][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_1  ( .A(\u_div/PartRem[19][1] ), .B(
        net32384), .CI(\u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[18][2] ), .S(
        \u_div/SumTmp[18][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_2  ( .A(\u_div/PartRem[19][2] ), .B(
        net32364), .CI(\u_div/CryTmp[18][2] ), .CO(\u_div/CryTmp[18][3] ), .S(
        \u_div/SumTmp[18][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_3  ( .A(\u_div/PartRem[19][3] ), .B(
        net32336), .CI(\u_div/CryTmp[18][3] ), .CO(\u_div/CryTmp[18][4] ), .S(
        \u_div/SumTmp[18][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_4  ( .A(\u_div/PartRem[19][4] ), .B(
        net32312), .CI(\u_div/CryTmp[18][4] ), .CO(\u_div/CryTmp[18][5] ), .S(
        \u_div/SumTmp[18][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_5  ( .A(\u_div/PartRem[19][5] ), .B(
        net32282), .CI(\u_div/CryTmp[18][5] ), .CO(\u_div/CryTmp[18][6] ), .S(
        \u_div/SumTmp[18][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_6  ( .A(\u_div/PartRem[19][6] ), .B(
        net32252), .CI(\u_div/CryTmp[18][6] ), .CO(\u_div/CryTmp[18][7] ), .S(
        \u_div/SumTmp[18][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_7  ( .A(\u_div/PartRem[19][7] ), .B(
        net32222), .CI(\u_div/CryTmp[18][7] ), .CO(\u_div/CryTmp[18][8] ), .S(
        \u_div/SumTmp[18][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_8  ( .A(\u_div/PartRem[19][8] ), .B(
        net32198), .CI(n137), .CO(\u_div/CryTmp[18][9] ), .S(
        \u_div/SumTmp[18][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_9  ( .A(\u_div/PartRem[19][9] ), .B(
        net32166), .CI(\u_div/CryTmp[18][9] ), .CO(\u_div/CryTmp[18][10] ), 
        .S(\u_div/SumTmp[18][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_10  ( .A(\u_div/PartRem[19][10] ), .B(
        net32142), .CI(\u_div/CryTmp[18][10] ), .CO(\u_div/CryTmp[18][11] ), 
        .S(\u_div/SumTmp[18][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_11  ( .A(\u_div/PartRem[19][11] ), .B(
        net32116), .CI(\u_div/CryTmp[18][11] ), .CO(\u_div/CryTmp[18][12] ), 
        .S(\u_div/SumTmp[18][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_12  ( .A(\u_div/PartRem[19][12] ), .B(
        net32090), .CI(\u_div/CryTmp[18][12] ), .CO(\u_div/CryTmp[18][13] ), 
        .S(\u_div/SumTmp[18][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_13  ( .A(\u_div/PartRem[19][13] ), .B(
        net32066), .CI(\u_div/CryTmp[18][13] ), .CO(\u_div/CryTmp[18][14] ), 
        .S(\u_div/SumTmp[18][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_14  ( .A(\u_div/PartRem[19][14] ), .B(
        net32044), .CI(\u_div/CryTmp[18][14] ), .CO(\u_div/CryTmp[18][15] ), 
        .S(\u_div/SumTmp[18][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_15  ( .A(\u_div/PartRem[19][15] ), .B(
        net32014), .CI(n626), .CO(\u_div/CryTmp[18][16] ), .S(
        \u_div/SumTmp[18][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_16  ( .A(\u_div/PartRem[19][16] ), .B(
        net31984), .CI(\u_div/CryTmp[18][16] ), .CO(\u_div/CryTmp[18][17] ), 
        .S(\u_div/SumTmp[18][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_17  ( .A(\u_div/CryTmp[18][17] ), .B(
        net31960), .CI(n633), .CO(\u_div/CryTmp[18][18] ), .S(
        \u_div/SumTmp[18][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_18  ( .A(\u_div/PartRem[19][18] ), .B(
        net31938), .CI(\u_div/CryTmp[18][18] ), .CO(\u_div/CryTmp[18][19] ), 
        .S(\u_div/SumTmp[18][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_19  ( .A(\u_div/PartRem[19][19] ), .B(
        net31912), .CI(\u_div/CryTmp[18][19] ), .CO(\u_div/CryTmp[18][20] ), 
        .S(\u_div/SumTmp[18][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_20  ( .A(\u_div/PartRem[19][20] ), .B(
        net31884), .CI(\u_div/CryTmp[18][20] ), .CO(\u_div/CryTmp[18][21] ), 
        .S(\u_div/SumTmp[18][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_21  ( .A(\u_div/PartRem[19][21] ), .B(
        net31856), .CI(\u_div/CryTmp[18][21] ), .CO(\u_div/CryTmp[18][22] ), 
        .S(\u_div/SumTmp[18][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_18_23  ( .A(\u_div/PartRem[19][23] ), .B(
        net31802), .CI(n133), .CO(\u_div/CryTmp[18][24] ), .S(
        \u_div/SumTmp[18][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_16_1  ( .A(\u_div/CryTmp[22][1] ), .B(
        net32384), .CI(\u_div/PartRem[17][1] ), .CO(\u_div/CryTmp[16][2] ), 
        .S(\u_div/SumTmp[16][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_21  ( .A(\u_div/PartRem[25][21] ), .B(
        net31854), .CI(n166), .CO(\u_div/CryTmp[24][22] ), .S(
        \u_div/SumTmp[24][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_1  ( .A(\u_div/PartRem[24][1] ), .B(
        net32384), .CI(\u_div/CryTmp[23][1] ), .CO(\u_div/CryTmp[23][2] ), .S(
        \u_div/SumTmp[23][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_2  ( .A(\u_div/PartRem[24][2] ), .B(
        net32364), .CI(\u_div/CryTmp[23][2] ), .CO(\u_div/CryTmp[23][3] ), .S(
        \u_div/SumTmp[23][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_3  ( .A(\u_div/PartRem[24][3] ), .B(
        net32336), .CI(\u_div/CryTmp[23][3] ), .CO(\u_div/CryTmp[23][4] ), .S(
        \u_div/SumTmp[23][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_4  ( .A(\u_div/PartRem[24][4] ), .B(
        net32312), .CI(\u_div/CryTmp[23][4] ), .CO(\u_div/CryTmp[23][5] ), .S(
        \u_div/SumTmp[23][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_5  ( .A(\u_div/PartRem[24][5] ), .B(
        net32282), .CI(\u_div/CryTmp[23][5] ), .CO(\u_div/CryTmp[23][6] ), .S(
        \u_div/SumTmp[23][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_6  ( .A(\u_div/PartRem[24][6] ), .B(
        net32252), .CI(\u_div/CryTmp[23][6] ), .CO(\u_div/CryTmp[23][7] ), .S(
        \u_div/SumTmp[23][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_7  ( .A(\u_div/PartRem[24][7] ), .B(
        net32222), .CI(\u_div/CryTmp[23][7] ), .CO(\u_div/CryTmp[23][8] ), .S(
        \u_div/SumTmp[23][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_8  ( .A(\u_div/PartRem[24][8] ), .B(
        net32198), .CI(n93), .CO(\u_div/CryTmp[23][9] ), .S(
        \u_div/SumTmp[23][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_9  ( .A(\u_div/PartRem[24][9] ), .B(
        net32166), .CI(\u_div/CryTmp[23][9] ), .CO(\u_div/CryTmp[23][10] ), 
        .S(\u_div/SumTmp[23][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_10  ( .A(\u_div/PartRem[24][10] ), .B(
        net32142), .CI(\u_div/CryTmp[23][10] ), .CO(\u_div/CryTmp[23][11] ), 
        .S(\u_div/SumTmp[23][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_11  ( .A(\u_div/PartRem[24][11] ), .B(
        net32116), .CI(\u_div/CryTmp[23][11] ), .CO(\u_div/CryTmp[23][12] ), 
        .S(\u_div/SumTmp[23][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_12  ( .A(\u_div/PartRem[24][12] ), .B(
        net32088), .CI(\u_div/CryTmp[23][12] ), .CO(\u_div/CryTmp[23][13] ), 
        .S(\u_div/SumTmp[23][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_13  ( .A(\u_div/PartRem[24][13] ), .B(
        net32078), .CI(\u_div/CryTmp[23][13] ), .CO(\u_div/CryTmp[23][14] ), 
        .S(\u_div/SumTmp[23][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_14  ( .A(\u_div/PartRem[24][14] ), .B(
        net32044), .CI(\u_div/CryTmp[23][14] ), .CO(\u_div/CryTmp[23][15] ), 
        .S(\u_div/SumTmp[23][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_15  ( .A(\u_div/PartRem[24][15] ), .B(
        net32014), .CI(\u_div/CryTmp[23][15] ), .CO(\u_div/CryTmp[23][16] ), 
        .S(\u_div/SumTmp[23][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_17  ( .A(\u_div/PartRem[24][17] ), .B(
        net31960), .CI(n567), .CO(\u_div/CryTmp[23][18] ), .S(
        \u_div/SumTmp[23][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_18  ( .A(\u_div/PartRem[24][18] ), .B(
        net31938), .CI(\u_div/CryTmp[23][18] ), .CO(\u_div/CryTmp[23][19] ), 
        .S(\u_div/SumTmp[23][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_19  ( .A(\u_div/PartRem[24][19] ), .B(
        net31912), .CI(\u_div/CryTmp[23][19] ), .CO(\u_div/CryTmp[23][20] ), 
        .S(\u_div/SumTmp[23][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_22  ( .A(\u_div/PartRem[24][22] ), .B(
        n135), .CI(net31828), .CO(\u_div/CryTmp[23][23] ), .S(
        \u_div/SumTmp[23][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_23  ( .A(n559), .B(net31802), .CI(
        \u_div/CryTmp[23][23] ), .CO(n1240), .S(\u_div/SumTmp[23][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_17  ( .A(\u_div/PartRem[23][17] ), .B(
        net31960), .CI(\u_div/CryTmp[22][17] ), .CO(\u_div/CryTmp[22][18] ), 
        .S(\u_div/SumTmp[22][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_18  ( .A(\u_div/PartRem[23][18] ), .B(
        net31938), .CI(n579), .CO(\u_div/CryTmp[22][19] ), .S(
        \u_div/SumTmp[22][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_19  ( .A(\u_div/PartRem[23][19] ), .B(
        net31912), .CI(\u_div/CryTmp[22][19] ), .CO(\u_div/CryTmp[22][20] ), 
        .S(\u_div/SumTmp[22][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_20  ( .A(\u_div/PartRem[23][20] ), .B(
        net31884), .CI(\u_div/CryTmp[22][20] ), .CO(\u_div/CryTmp[22][21] ), 
        .S(\u_div/SumTmp[22][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_21  ( .A(\u_div/PartRem[23][21] ), .B(
        net31856), .CI(\u_div/CryTmp[22][21] ), .CO(\u_div/CryTmp[22][22] ), 
        .S(\u_div/SumTmp[22][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_22  ( .A(\u_div/PartRem[23][22] ), .B(
        net31828), .CI(\u_div/CryTmp[22][22] ), .CO(\u_div/CryTmp[22][23] ), 
        .S(\u_div/SumTmp[22][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_23  ( .A(\u_div/PartRem[23][23] ), .B(
        n577), .CI(net31802), .CO(\u_div/CryTmp[22][24] ), .S(
        \u_div/SumTmp[22][23] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_1  ( .A(\u_div/PartRem[23][1] ), .B(
        net32384), .CI(\u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[22][2] ), .S(
        \u_div/SumTmp[22][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_2  ( .A(\u_div/PartRem[23][2] ), .B(
        net32364), .CI(\u_div/CryTmp[22][2] ), .CO(\u_div/CryTmp[22][3] ), .S(
        \u_div/SumTmp[22][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_3  ( .A(\u_div/PartRem[23][3] ), .B(
        net32336), .CI(\u_div/CryTmp[22][3] ), .CO(\u_div/CryTmp[22][4] ), .S(
        \u_div/SumTmp[22][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_4  ( .A(\u_div/PartRem[23][4] ), .B(
        net32312), .CI(\u_div/CryTmp[22][4] ), .CO(\u_div/CryTmp[22][5] ), .S(
        \u_div/SumTmp[22][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_22_5  ( .A(\u_div/PartRem[23][5] ), .B(
        net32282), .CI(\u_div/CryTmp[22][5] ), .CO(\u_div/CryTmp[22][6] ), .S(
        \u_div/SumTmp[22][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_1  ( .A(\u_div/PartRem[22][1] ), .B(
        net32384), .CI(\u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[21][2] ), .S(
        \u_div/SumTmp[21][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_2  ( .A(\u_div/PartRem[22][2] ), .B(
        net32364), .CI(\u_div/CryTmp[21][2] ), .CO(\u_div/CryTmp[21][3] ), .S(
        \u_div/SumTmp[21][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_3  ( .A(\u_div/PartRem[22][3] ), .B(
        net32336), .CI(\u_div/CryTmp[21][3] ), .CO(\u_div/CryTmp[21][4] ), .S(
        \u_div/SumTmp[21][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_5  ( .A(n562), .B(net32282), .CI(
        net46688), .CO(\u_div/CryTmp[21][6] ), .S(\u_div/SumTmp[21][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_7  ( .A(\u_div/PartRem[22][7] ), .B(
        net32222), .CI(n314), .CO(\u_div/CryTmp[21][8] ), .S(
        \u_div/SumTmp[21][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_8  ( .A(\u_div/PartRem[22][8] ), .B(
        net32198), .CI(\u_div/CryTmp[21][8] ), .CO(\u_div/CryTmp[21][9] ), .S(
        \u_div/SumTmp[21][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_9  ( .A(\u_div/PartRem[22][9] ), .B(
        net32166), .CI(n182), .CO(\u_div/CryTmp[21][10] ), .S(
        \u_div/SumTmp[21][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_10  ( .A(\u_div/PartRem[22][10] ), .B(
        net32142), .CI(\u_div/CryTmp[21][10] ), .CO(\u_div/CryTmp[21][11] ), 
        .S(\u_div/SumTmp[21][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_11  ( .A(\u_div/PartRem[22][11] ), .B(
        net32116), .CI(\u_div/CryTmp[21][11] ), .CO(\u_div/CryTmp[21][12] ), 
        .S(\u_div/SumTmp[21][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_17  ( .A(\u_div/PartRem[21][17] ), .B(
        net31960), .CI(n111), .CO(\u_div/CryTmp[20][18] ), .S(
        \u_div/SumTmp[20][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_1  ( .A(n565), .B(net32384), .CI(
        \u_div/CryTmp[22][1] ), .CO(\u_div/CryTmp[20][2] ), .S(
        \u_div/SumTmp[20][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_2  ( .A(\u_div/PartRem[21][2] ), .B(
        net32364), .CI(\u_div/CryTmp[20][2] ), .CO(\u_div/CryTmp[20][3] ), .S(
        \u_div/SumTmp[20][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_3  ( .A(\u_div/PartRem[21][3] ), .B(
        net32336), .CI(\u_div/CryTmp[20][3] ), .CO(\u_div/CryTmp[20][4] ), .S(
        \u_div/SumTmp[20][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_4  ( .A(\u_div/PartRem[21][4] ), .B(
        net32312), .CI(\u_div/CryTmp[20][4] ), .CO(\u_div/CryTmp[20][5] ), .S(
        \u_div/SumTmp[20][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_5  ( .A(\u_div/PartRem[21][5] ), .B(
        net32282), .CI(\u_div/CryTmp[20][5] ), .CO(\u_div/CryTmp[20][6] ), .S(
        \u_div/SumTmp[20][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_6  ( .A(\u_div/PartRem[21][6] ), .B(
        net32252), .CI(n571), .CO(\u_div/CryTmp[20][7] ), .S(
        \u_div/SumTmp[20][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_7  ( .A(\u_div/PartRem[21][7] ), .B(
        net32222), .CI(\u_div/CryTmp[20][7] ), .CO(\u_div/CryTmp[20][8] ), .S(
        \u_div/SumTmp[20][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_8  ( .A(n581), .B(net32198), .CI(n572), 
        .CO(\u_div/CryTmp[20][9] ), .S(\u_div/SumTmp[20][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_9  ( .A(\u_div/PartRem[21][9] ), .B(
        net32166), .CI(\u_div/CryTmp[20][9] ), .CO(\u_div/CryTmp[20][10] ), 
        .S(\u_div/SumTmp[20][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_10  ( .A(\u_div/PartRem[21][10] ), .B(
        net32142), .CI(\u_div/CryTmp[20][10] ), .CO(\u_div/CryTmp[20][11] ), 
        .S(\u_div/SumTmp[20][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_11  ( .A(\u_div/PartRem[21][11] ), .B(
        net32116), .CI(n246), .CO(\u_div/CryTmp[20][12] ), .S(
        \u_div/SumTmp[20][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_13  ( .A(\u_div/PartRem[21][13] ), .B(
        net32066), .CI(n85), .CO(\u_div/CryTmp[20][14] ), .S(
        \u_div/SumTmp[20][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_15  ( .A(\u_div/PartRem[21][15] ), .B(
        net32014), .CI(n175), .CO(\u_div/CryTmp[20][16] ), .S(
        \u_div/SumTmp[20][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_20_16  ( .A(\u_div/PartRem[21][16] ), .B(
        net31982), .CI(\u_div/CryTmp[20][16] ), .CO(\u_div/CryTmp[20][17] ), 
        .S(\u_div/SumTmp[20][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_18  ( .A(\u_div/PartRem[20][18] ), .B(
        net31938), .CI(\u_div/CryTmp[19][18] ), .CO(\u_div/CryTmp[19][19] ), 
        .S(\u_div/SumTmp[19][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_1  ( .A(net32384), .B(
        \u_div/PartRem[20][1] ), .CI(\u_div/CryTmp[22][1] ), .CO(
        \u_div/CryTmp[19][2] ), .S(\u_div/SumTmp[19][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_2  ( .A(\u_div/PartRem[20][2] ), .B(
        net32364), .CI(\u_div/CryTmp[19][2] ), .CO(\u_div/CryTmp[19][3] ), .S(
        \u_div/SumTmp[19][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_3  ( .A(\u_div/PartRem[20][3] ), .B(
        net32336), .CI(\u_div/CryTmp[19][3] ), .CO(\u_div/CryTmp[19][4] ), .S(
        \u_div/SumTmp[19][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_4  ( .A(\u_div/PartRem[20][4] ), .B(
        net32312), .CI(\u_div/CryTmp[19][4] ), .CO(\u_div/CryTmp[19][5] ), .S(
        \u_div/SumTmp[19][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_5  ( .A(\u_div/PartRem[20][5] ), .B(
        net32282), .CI(\u_div/CryTmp[19][5] ), .CO(\u_div/CryTmp[19][6] ), .S(
        \u_div/SumTmp[19][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_6  ( .A(\u_div/PartRem[20][6] ), .B(
        net32252), .CI(\u_div/CryTmp[19][6] ), .CO(\u_div/CryTmp[19][7] ), .S(
        \u_div/SumTmp[19][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_7  ( .A(\u_div/PartRem[20][7] ), .B(
        net32222), .CI(\u_div/CryTmp[19][7] ), .CO(\u_div/CryTmp[19][8] ), .S(
        \u_div/SumTmp[19][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_8  ( .A(\u_div/PartRem[20][8] ), .B(
        net32198), .CI(\u_div/CryTmp[19][8] ), .CO(\u_div/CryTmp[19][9] ), .S(
        \u_div/SumTmp[19][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_10  ( .A(\u_div/PartRem[20][10] ), .B(
        n564), .CI(net32142), .CO(\u_div/CryTmp[19][11] ), .S(
        \u_div/SumTmp[19][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_11  ( .A(\u_div/PartRem[20][11] ), .B(
        net32116), .CI(\u_div/CryTmp[19][11] ), .CO(\u_div/CryTmp[19][12] ), 
        .S(\u_div/SumTmp[19][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_12  ( .A(\u_div/PartRem[20][12] ), .B(
        net32090), .CI(\u_div/CryTmp[19][12] ), .CO(\u_div/CryTmp[19][13] ), 
        .S(\u_div/SumTmp[19][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_14  ( .A(n588), .B(net32044), .CI(n575), 
        .CO(\u_div/CryTmp[19][15] ), .S(\u_div/SumTmp[19][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_15  ( .A(n586), .B(net32014), .CI(
        \u_div/CryTmp[19][15] ), .CO(\u_div/CryTmp[19][16] ), .S(
        \u_div/SumTmp[19][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_16  ( .A(n590), .B(net31982), .CI(
        \u_div/CryTmp[19][16] ), .CO(\u_div/CryTmp[19][17] ), .S(
        \u_div/SumTmp[19][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_17  ( .A(\u_div/PartRem[20][17] ), .B(
        net31960), .CI(\u_div/CryTmp[19][17] ), .CO(\u_div/CryTmp[19][18] ), 
        .S(\u_div/SumTmp[19][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_14  ( .A(\u_div/PartRem[26][14] ), .B(
        net32046), .CI(\u_div/CryTmp[25][14] ), .CO(\u_div/CryTmp[25][15] ), 
        .S(\u_div/SumTmp[25][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_15  ( .A(\u_div/PartRem[26][15] ), .B(
        net32016), .CI(\u_div/CryTmp[25][15] ), .CO(\u_div/CryTmp[25][16] ), 
        .S(\u_div/SumTmp[25][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_16  ( .A(\u_div/PartRem[26][16] ), .B(
        net31982), .CI(\u_div/CryTmp[25][16] ), .CO(\u_div/CryTmp[25][17] ), 
        .S(\u_div/SumTmp[25][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_17  ( .A(\u_div/PartRem[26][17] ), .B(
        net31960), .CI(\u_div/CryTmp[25][17] ), .CO(\u_div/CryTmp[25][18] ), 
        .S(\u_div/SumTmp[25][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_19  ( .A(\u_div/PartRem[26][19] ), .B(
        net31914), .CI(n292), .CO(\u_div/CryTmp[25][20] ), .S(
        \u_div/SumTmp[25][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_20  ( .A(\u_div/PartRem[26][20] ), .B(
        net31884), .CI(\u_div/CryTmp[25][20] ), .CO(\u_div/CryTmp[25][21] ), 
        .S(\u_div/SumTmp[25][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_1  ( .A(\u_div/PartRem[26][1] ), .B(
        net32386), .CI(\u_div/CryTmp[25][1] ), .CO(\u_div/CryTmp[25][2] ), .S(
        \u_div/SumTmp[25][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_2  ( .A(\u_div/PartRem[26][2] ), .B(
        net32366), .CI(\u_div/CryTmp[25][2] ), .CO(\u_div/CryTmp[25][3] ), .S(
        \u_div/SumTmp[25][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_3  ( .A(\u_div/PartRem[26][3] ), .B(
        net32338), .CI(\u_div/CryTmp[25][3] ), .CO(\u_div/CryTmp[25][4] ), .S(
        \u_div/SumTmp[25][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_4  ( .A(\u_div/PartRem[26][4] ), .B(n504), .CI(net32314), .CO(\u_div/CryTmp[25][5] ), .S(\u_div/SumTmp[25][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_5  ( .A(\u_div/PartRem[26][5] ), .B(
        net32284), .CI(\u_div/CryTmp[25][5] ), .CO(\u_div/CryTmp[25][6] ), .S(
        \u_div/SumTmp[25][5] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_25_6  ( .A(\u_div/PartRem[26][6] ), .B(
        net32254), .CI(\u_div/CryTmp[25][6] ), .CO(\u_div/CryTmp[25][7] ), .S(
        \u_div/SumTmp[25][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_7  ( .A(\u_div/PartRem[26][7] ), .B(
        net32222), .CI(n512), .CO(\u_div/CryTmp[25][8] ), .S(
        \u_div/SumTmp[25][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_8  ( .A(net32200), .B(
        \u_div/CryTmp[25][8] ), .CI(\u_div/PartRem[26][8] ), .CO(
        \u_div/CryTmp[25][9] ), .S(\u_div/SumTmp[25][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_9  ( .A(\u_div/PartRem[26][9] ), .B(
        net32166), .CI(n521), .CO(\u_div/CryTmp[25][10] ), .S(
        \u_div/SumTmp[25][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_11  ( .A(\u_div/PartRem[26][11] ), .B(
        net49055), .CI(n322), .CO(\u_div/CryTmp[25][12] ), .S(
        \u_div/SumTmp[25][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_12  ( .A(\u_div/PartRem[26][12] ), .B(
        net32088), .CI(\u_div/CryTmp[25][12] ), .CO(\u_div/CryTmp[25][13] ), 
        .S(\u_div/SumTmp[25][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_13  ( .A(\u_div/PartRem[26][13] ), .B(
        n519), .CI(net32078), .CO(\u_div/CryTmp[25][14] ), .S(
        \u_div/SumTmp[25][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_20  ( .A(\u_div/PartRem[25][20] ), .B(
        net31884), .CI(\u_div/CryTmp[24][20] ), .CO(\u_div/CryTmp[24][21] ), 
        .S(\u_div/SumTmp[24][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_2  ( .A(\u_div/PartRem[25][2] ), .B(
        net32366), .CI(\u_div/CryTmp[24][2] ), .CO(\u_div/CryTmp[24][3] ), .S(
        \u_div/SumTmp[24][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_3  ( .A(\u_div/PartRem[25][3] ), .B(
        net32338), .CI(\u_div/CryTmp[24][3] ), .CO(\u_div/CryTmp[24][4] ), .S(
        \u_div/SumTmp[24][3] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_24_4  ( .A(\u_div/PartRem[25][4] ), .B(
        net32314), .CI(\u_div/CryTmp[24][4] ), .CO(\u_div/CryTmp[24][5] ), .S(
        \u_div/SumTmp[24][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_5  ( .A(\u_div/PartRem[25][5] ), .B(
        net32284), .CI(n508), .CO(\u_div/CryTmp[24][6] ), .S(
        \u_div/SumTmp[24][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_6  ( .A(\u_div/PartRem[25][6] ), .B(
        net32254), .CI(\u_div/CryTmp[24][6] ), .CO(\u_div/CryTmp[24][7] ), .S(
        \u_div/SumTmp[24][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_7  ( .A(\u_div/PartRem[25][7] ), .B(
        net32222), .CI(\u_div/CryTmp[24][7] ), .CO(\u_div/CryTmp[24][8] ), .S(
        \u_div/SumTmp[24][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_8  ( .A(\u_div/PartRem[25][8] ), .B(
        net32200), .CI(\u_div/CryTmp[24][8] ), .CO(\u_div/CryTmp[24][9] ), .S(
        \u_div/SumTmp[24][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_9  ( .A(n180), .B(net32166), .CI(
        \u_div/CryTmp[24][9] ), .CO(\u_div/CryTmp[24][10] ), .S(
        \u_div/SumTmp[24][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_10  ( .A(\u_div/PartRem[25][10] ), .B(
        net32140), .CI(n510), .CO(\u_div/CryTmp[24][11] ), .S(
        \u_div/SumTmp[24][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_11  ( .A(\u_div/PartRem[25][11] ), .B(
        net49055), .CI(\u_div/CryTmp[24][11] ), .CO(\u_div/CryTmp[24][12] ), 
        .S(\u_div/SumTmp[24][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_12  ( .A(\u_div/PartRem[25][12] ), .B(
        net32088), .CI(\u_div/CryTmp[24][12] ), .CO(\u_div/CryTmp[24][13] ), 
        .S(\u_div/SumTmp[24][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_13  ( .A(\u_div/PartRem[25][13] ), .B(
        net32078), .CI(n514), .CO(\u_div/CryTmp[24][14] ), .S(
        \u_div/SumTmp[24][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_14  ( .A(\u_div/PartRem[25][14] ), .B(
        net32046), .CI(n516), .CO(\u_div/CryTmp[24][15] ), .S(
        \u_div/SumTmp[24][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_15  ( .A(\u_div/PartRem[25][15] ), .B(
        net32016), .CI(\u_div/CryTmp[24][15] ), .CO(\u_div/CryTmp[24][16] ), 
        .S(\u_div/SumTmp[24][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_16  ( .A(\u_div/PartRem[25][16] ), .B(
        net31982), .CI(\u_div/CryTmp[24][16] ), .CO(\u_div/CryTmp[24][17] ), 
        .S(\u_div/SumTmp[24][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_17  ( .A(\u_div/PartRem[25][17] ), .B(
        net31960), .CI(\u_div/CryTmp[24][17] ), .CO(\u_div/CryTmp[24][18] ), 
        .S(\u_div/SumTmp[24][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_18  ( .A(\u_div/PartRem[25][18] ), .B(
        net31938), .CI(\u_div/CryTmp[24][18] ), .CO(\u_div/CryTmp[24][19] ), 
        .S(\u_div/SumTmp[24][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_19  ( .A(\u_div/PartRem[25][19] ), .B(
        net31914), .CI(\u_div/CryTmp[24][19] ), .CO(\u_div/CryTmp[24][20] ), 
        .S(\u_div/SumTmp[24][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_1  ( .A(\u_div/PartRem[30][1] ), .B(
        net32386), .CI(\u_div/CryTmp[29][1] ), .CO(\u_div/CryTmp[29][2] ), .S(
        \u_div/SumTmp[29][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_2  ( .A(\u_div/PartRem[30][2] ), .B(
        net32366), .CI(\u_div/CryTmp[29][2] ), .CO(\u_div/CryTmp[29][3] ), .S(
        \u_div/SumTmp[29][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_3  ( .A(\u_div/PartRem[30][3] ), .B(
        net32338), .CI(\u_div/CryTmp[29][3] ), .CO(\u_div/CryTmp[29][4] ), .S(
        \u_div/SumTmp[29][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_4  ( .A(\u_div/PartRem[30][4] ), .B(
        net32314), .CI(\u_div/CryTmp[29][4] ), .CO(\u_div/CryTmp[29][5] ), .S(
        \u_div/SumTmp[29][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_5  ( .A(\u_div/PartRem[30][5] ), .B(
        net32284), .CI(\u_div/CryTmp[29][5] ), .CO(\u_div/CryTmp[29][6] ), .S(
        \u_div/SumTmp[29][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_6  ( .A(\u_div/PartRem[30][6] ), .B(
        net32254), .CI(\u_div/CryTmp[29][6] ), .CO(\u_div/CryTmp[29][7] ), .S(
        \u_div/SumTmp[29][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_7  ( .A(\u_div/PartRem[30][7] ), .B(
        net32222), .CI(\u_div/CryTmp[29][7] ), .CO(\u_div/CryTmp[29][8] ), .S(
        \u_div/SumTmp[29][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_8  ( .A(\u_div/PartRem[30][8] ), .B(
        net32200), .CI(\u_div/CryTmp[29][8] ), .CO(\u_div/CryTmp[29][9] ), .S(
        \u_div/SumTmp[29][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_10  ( .A(\u_div/PartRem[30][10] ), .B(
        net32140), .CI(n248), .CO(\u_div/CryTmp[29][11] ), .S(
        \u_div/SumTmp[29][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_11  ( .A(\u_div/PartRem[30][11] ), .B(
        net49055), .CI(\u_div/CryTmp[29][11] ), .CO(\u_div/CryTmp[29][12] ), 
        .S(\u_div/SumTmp[29][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_12  ( .A(\u_div/PartRem[30][12] ), .B(
        net32088), .CI(\u_div/CryTmp[29][12] ), .CO(\u_div/CryTmp[29][13] ), 
        .S(\u_div/SumTmp[29][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_13  ( .A(\u_div/PartRem[30][13] ), .B(
        net32078), .CI(\u_div/CryTmp[29][13] ), .CO(\u_div/CryTmp[29][14] ), 
        .S(\u_div/SumTmp[29][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_14  ( .A(\u_div/PartRem[30][14] ), .B(
        net32046), .CI(\u_div/CryTmp[29][14] ), .CO(\u_div/CryTmp[29][15] ), 
        .S(\u_div/SumTmp[29][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_15  ( .A(\u_div/PartRem[30][15] ), .B(
        net32016), .CI(\u_div/CryTmp[29][15] ), .CO(\u_div/CryTmp[29][16] ), 
        .S(\u_div/SumTmp[29][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_16  ( .A(\u_div/PartRem[30][16] ), .B(
        net31982), .CI(n498), .CO(\u_div/CryTmp[29][17] ), .S(
        \u_div/SumTmp[29][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_29_17  ( .A(\u_div/PartRem[30][17] ), .B(
        net31960), .CI(\u_div/CryTmp[29][17] ), .CO(\u_div/CryTmp[29][18] ), 
        .S(\u_div/SumTmp[29][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_1  ( .A(\u_div/CryTmp[28][1] ), .B(
        net32386), .CI(\u_div/PartRem[29][1] ), .CO(\u_div/CryTmp[28][2] ), 
        .S(\u_div/SumTmp[28][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_2  ( .A(\u_div/PartRem[29][2] ), .B(
        net32366), .CI(\u_div/CryTmp[28][2] ), .CO(\u_div/CryTmp[28][3] ), .S(
        \u_div/SumTmp[28][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_3  ( .A(\u_div/PartRem[29][3] ), .B(
        net32338), .CI(\u_div/CryTmp[28][3] ), .CO(\u_div/CryTmp[28][4] ), .S(
        \u_div/SumTmp[28][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_4  ( .A(\u_div/PartRem[29][4] ), .B(
        net32314), .CI(\u_div/CryTmp[28][4] ), .CO(\u_div/CryTmp[28][5] ), .S(
        \u_div/SumTmp[28][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_5  ( .A(\u_div/PartRem[29][5] ), .B(
        net32284), .CI(\u_div/CryTmp[28][5] ), .CO(\u_div/CryTmp[28][6] ), .S(
        \u_div/SumTmp[28][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_6  ( .A(\u_div/PartRem[29][6] ), .B(
        net32254), .CI(\u_div/CryTmp[28][6] ), .CO(\u_div/CryTmp[28][7] ), .S(
        \u_div/SumTmp[28][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_7  ( .A(\u_div/PartRem[29][7] ), .B(
        net32224), .CI(\u_div/CryTmp[28][7] ), .CO(\u_div/CryTmp[28][8] ), .S(
        \u_div/SumTmp[28][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_8  ( .A(\u_div/PartRem[29][8] ), .B(
        net32200), .CI(\u_div/CryTmp[28][8] ), .CO(\u_div/CryTmp[28][9] ), .S(
        \u_div/SumTmp[28][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_28_9  ( .A(\u_div/PartRem[29][9] ), .B(
        net32166), .CI(\u_div/CryTmp[28][9] ), .CO(\u_div/CryTmp[28][10] ), 
        .S(\u_div/SumTmp[28][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_1  ( .A(\u_div/PartRem[28][1] ), .B(
        net32386), .CI(\u_div/CryTmp[27][1] ), .CO(\u_div/CryTmp[27][2] ), .S(
        \u_div/SumTmp[27][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_2  ( .A(\u_div/PartRem[28][2] ), .B(
        net32366), .CI(\u_div/CryTmp[27][2] ), .CO(\u_div/CryTmp[27][3] ), .S(
        \u_div/SumTmp[27][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_3  ( .A(\u_div/PartRem[28][3] ), .B(
        net32338), .CI(n488), .CO(\u_div/CryTmp[27][4] ), .S(
        \u_div/SumTmp[27][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_4  ( .A(\u_div/PartRem[28][4] ), .B(
        net32314), .CI(\u_div/CryTmp[27][4] ), .CO(\u_div/CryTmp[27][5] ), .S(
        \u_div/SumTmp[27][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_5  ( .A(\u_div/PartRem[28][5] ), .B(
        net32284), .CI(\u_div/CryTmp[27][5] ), .CO(\u_div/CryTmp[27][6] ), .S(
        \u_div/SumTmp[27][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_6  ( .A(\u_div/PartRem[28][6] ), .B(
        net32254), .CI(\u_div/CryTmp[27][6] ), .CO(\u_div/CryTmp[27][7] ), .S(
        \u_div/SumTmp[27][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_7  ( .A(\u_div/PartRem[28][7] ), .B(
        net32222), .CI(\u_div/CryTmp[27][7] ), .CO(\u_div/CryTmp[27][8] ), .S(
        \u_div/SumTmp[27][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_9  ( .A(\u_div/PartRem[28][9] ), .B(
        net32168), .CI(n236), .CO(\u_div/CryTmp[27][10] ), .S(
        \u_div/SumTmp[27][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_27_10  ( .A(\u_div/PartRem[28][10] ), .B(
        net32142), .CI(\u_div/CryTmp[27][10] ), .CO(\u_div/CryTmp[27][11] ), 
        .S(\u_div/SumTmp[27][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_1  ( .A(\u_div/PartRem[27][1] ), .B(
        net32386), .CI(\u_div/CryTmp[26][1] ), .CO(\u_div/CryTmp[26][2] ), .S(
        \u_div/SumTmp[26][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_2  ( .A(\u_div/PartRem[27][2] ), .B(
        net32366), .CI(\u_div/CryTmp[26][2] ), .CO(\u_div/CryTmp[26][3] ), .S(
        \u_div/SumTmp[26][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_4  ( .A(\u_div/PartRem[27][4] ), .B(
        net32314), .CI(n492), .CO(\u_div/CryTmp[26][5] ), .S(
        \u_div/SumTmp[26][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_5  ( .A(\u_div/CryTmp[26][5] ), .B(
        net32284), .CI(\u_div/PartRem[27][5] ), .CO(\u_div/CryTmp[26][6] ), 
        .S(\u_div/SumTmp[26][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_6  ( .A(\u_div/PartRem[27][6] ), .B(
        net32254), .CI(\u_div/CryTmp[26][6] ), .CO(\u_div/CryTmp[26][7] ), .S(
        \u_div/SumTmp[26][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_8  ( .A(\u_div/PartRem[27][8] ), .B(
        net32200), .CI(\u_div/CryTmp[26][8] ), .CO(\u_div/CryTmp[26][9] ), .S(
        \u_div/SumTmp[26][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_10  ( .A(net32140), .B(
        \u_div/PartRem[27][10] ), .CI(n250), .CO(\u_div/CryTmp[26][11] ), .S(
        \u_div/SumTmp[26][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_11  ( .A(n494), .B(net49055), .CI(
        \u_div/PartRem[27][11] ), .CO(\u_div/CryTmp[26][12] ), .S(
        \u_div/SumTmp[26][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_12  ( .A(\u_div/CryTmp[26][12] ), .B(
        net32088), .CI(\u_div/PartRem[27][12] ), .CO(\u_div/CryTmp[26][13] ), 
        .S(\u_div/SumTmp[26][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_13  ( .A(n28), .B(net32078), .CI(n178), 
        .CO(\u_div/CryTmp[26][14] ), .S(\u_div/SumTmp[26][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_14  ( .A(\u_div/PartRem[27][14] ), .B(
        net32046), .CI(\u_div/CryTmp[26][14] ), .CO(\u_div/CryTmp[26][15] ), 
        .S(\u_div/SumTmp[26][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_15  ( .A(\u_div/PartRem[27][15] ), .B(
        net32016), .CI(\u_div/CryTmp[26][15] ), .CO(\u_div/CryTmp[26][16] ), 
        .S(\u_div/SumTmp[26][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_16  ( .A(\u_div/PartRem[27][16] ), .B(
        net31982), .CI(\u_div/CryTmp[26][16] ), .CO(\u_div/CryTmp[26][17] ), 
        .S(\u_div/SumTmp[26][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_17  ( .A(\u_div/PartRem[27][17] ), .B(
        net31960), .CI(\u_div/CryTmp[26][17] ), .CO(\u_div/CryTmp[26][18] ), 
        .S(\u_div/SumTmp[26][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_18  ( .A(\u_div/PartRem[27][18] ), .B(
        net31938), .CI(\u_div/CryTmp[26][18] ), .CO(\u_div/CryTmp[26][19] ), 
        .S(\u_div/SumTmp[26][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_19  ( .A(\u_div/PartRem[27][19] ), .B(
        net31914), .CI(\u_div/CryTmp[26][19] ), .CO(\u_div/CryTmp[26][20] ), 
        .S(\u_div/SumTmp[26][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_20  ( .A(\u_div/PartRem[27][20] ), .B(
        net31882), .CI(\u_div/CryTmp[26][20] ), .CO(\u_div/CryTmp[26][21] ), 
        .S(\u_div/SumTmp[26][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_1  ( .A(\u_div/PartRem[37][1] ), .B(
        net32382), .CI(\u_div/CryTmp[36][1] ), .CO(\u_div/CryTmp[36][2] ), .S(
        \u_div/SumTmp[36][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_2  ( .A(\u_div/PartRem[37][2] ), .B(
        net32368), .CI(\u_div/CryTmp[36][2] ), .CO(\u_div/CryTmp[36][3] ), .S(
        \u_div/SumTmp[36][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_3  ( .A(\u_div/PartRem[37][3] ), .B(
        net32354), .CI(\u_div/CryTmp[36][3] ), .CO(\u_div/CryTmp[36][4] ), .S(
        \u_div/SumTmp[36][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_1  ( .A(\u_div/PartRem[36][1] ), .B(
        net32386), .CI(\u_div/CryTmp[35][1] ), .CO(\u_div/CryTmp[35][2] ), .S(
        \u_div/SumTmp[35][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_2  ( .A(\u_div/PartRem[36][2] ), .B(
        net32366), .CI(\u_div/CryTmp[35][2] ), .CO(\u_div/CryTmp[35][3] ), .S(
        \u_div/SumTmp[35][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_3  ( .A(\u_div/PartRem[36][3] ), .B(
        net32338), .CI(\u_div/CryTmp[35][3] ), .CO(\u_div/CryTmp[35][4] ), .S(
        \u_div/SumTmp[35][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_4  ( .A(\u_div/PartRem[36][4] ), .B(
        net32314), .CI(\u_div/CryTmp[35][4] ), .CO(\u_div/CryTmp[35][5] ), .S(
        \u_div/SumTmp[35][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_1  ( .A(n234), .B(net32386), .CI(
        \u_div/CryTmp[34][1] ), .CO(\u_div/CryTmp[34][2] ), .S(
        \u_div/SumTmp[34][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_2  ( .A(\u_div/PartRem[35][2] ), .B(
        net32366), .CI(\u_div/CryTmp[34][2] ), .CO(\u_div/CryTmp[34][3] ), .S(
        \u_div/SumTmp[34][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_3  ( .A(\u_div/PartRem[35][3] ), .B(
        net32338), .CI(\u_div/CryTmp[34][3] ), .CO(\u_div/CryTmp[34][4] ), .S(
        \u_div/SumTmp[34][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_4  ( .A(\u_div/PartRem[35][4] ), .B(
        net32314), .CI(\u_div/CryTmp[34][4] ), .CO(\u_div/CryTmp[34][5] ), .S(
        \u_div/SumTmp[34][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_5  ( .A(\u_div/PartRem[35][5] ), .B(
        net32284), .CI(\u_div/CryTmp[34][5] ), .CO(\u_div/CryTmp[34][6] ), .S(
        \u_div/SumTmp[34][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_6  ( .A(\u_div/PartRem[35][6] ), .B(
        net32254), .CI(\u_div/CryTmp[34][6] ), .CO(\u_div/CryTmp[34][7] ), .S(
        \u_div/SumTmp[34][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_7  ( .A(\u_div/PartRem[35][7] ), .B(
        net32242), .CI(\u_div/CryTmp[34][7] ), .CO(\u_div/CryTmp[34][8] ), .S(
        \u_div/SumTmp[34][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_9  ( .A(\u_div/PartRem[35][9] ), .B(
        net32186), .CI(\u_div/CryTmp[34][9] ), .CO(\u_div/CryTmp[34][10] ), 
        .S(\u_div/SumTmp[34][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_1  ( .A(\u_div/PartRem[34][1] ), .B(
        net32386), .CI(\u_div/CryTmp[33][1] ), .CO(\u_div/CryTmp[33][2] ), .S(
        \u_div/SumTmp[33][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_2  ( .A(\u_div/PartRem[34][2] ), .B(
        net32366), .CI(\u_div/CryTmp[33][2] ), .CO(\u_div/CryTmp[33][3] ), .S(
        \u_div/SumTmp[33][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_3  ( .A(\u_div/PartRem[34][3] ), .B(
        net32338), .CI(\u_div/CryTmp[33][3] ), .CO(\u_div/CryTmp[33][4] ), .S(
        \u_div/SumTmp[33][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_4  ( .A(\u_div/PartRem[34][4] ), .B(
        net32314), .CI(\u_div/CryTmp[33][4] ), .CO(\u_div/CryTmp[33][5] ), .S(
        \u_div/SumTmp[33][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_5  ( .A(\u_div/PartRem[34][5] ), .B(
        net32284), .CI(\u_div/CryTmp[33][5] ), .CO(\u_div/CryTmp[33][6] ), .S(
        \u_div/SumTmp[33][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_6  ( .A(\u_div/PartRem[34][6] ), .B(
        net32254), .CI(\u_div/CryTmp[33][6] ), .CO(\u_div/CryTmp[33][7] ), .S(
        \u_div/SumTmp[33][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_7  ( .A(\u_div/PartRem[34][7] ), .B(
        net32226), .CI(\u_div/CryTmp[33][7] ), .CO(\u_div/CryTmp[33][8] ), .S(
        \u_div/SumTmp[33][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_8  ( .A(\u_div/PartRem[34][8] ), .B(
        net32200), .CI(\u_div/CryTmp[33][8] ), .CO(\u_div/CryTmp[33][9] ), .S(
        \u_div/SumTmp[33][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_9  ( .A(\u_div/PartRem[34][9] ), .B(
        net32186), .CI(\u_div/CryTmp[33][9] ), .CO(\u_div/CryTmp[33][10] ), 
        .S(\u_div/SumTmp[33][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_33_10  ( .A(\u_div/CryTmp[33][10] ), .B(
        net32140), .CI(\u_div/PartRem[34][10] ), .CO(\u_div/CryTmp[33][11] ), 
        .S(\u_div/SumTmp[33][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_14  ( .A(\u_div/PartRem[33][14] ), .B(
        net32046), .CI(\u_div/CryTmp[32][14] ), .CO(\u_div/CryTmp[32][15] ), 
        .S(\u_div/SumTmp[32][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_1  ( .A(\u_div/PartRem[33][1] ), .B(
        net32386), .CI(\u_div/CryTmp[32][1] ), .CO(\u_div/CryTmp[32][2] ), .S(
        \u_div/SumTmp[32][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_2  ( .A(\u_div/PartRem[33][2] ), .B(
        net32366), .CI(\u_div/CryTmp[32][2] ), .CO(\u_div/CryTmp[32][3] ), .S(
        \u_div/SumTmp[32][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_3  ( .A(\u_div/PartRem[33][3] ), .B(
        net32338), .CI(\u_div/CryTmp[32][3] ), .CO(\u_div/CryTmp[32][4] ), .S(
        \u_div/SumTmp[32][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_4  ( .A(\u_div/PartRem[33][4] ), .B(
        net32314), .CI(\u_div/CryTmp[32][4] ), .CO(\u_div/CryTmp[32][5] ), .S(
        \u_div/SumTmp[32][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_5  ( .A(\u_div/PartRem[33][5] ), .B(
        net32284), .CI(\u_div/CryTmp[32][5] ), .CO(\u_div/CryTmp[32][6] ), .S(
        \u_div/SumTmp[32][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_6  ( .A(\u_div/PartRem[33][6] ), .B(
        net32254), .CI(\u_div/CryTmp[32][6] ), .CO(\u_div/CryTmp[32][7] ), .S(
        \u_div/SumTmp[32][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_7  ( .A(\u_div/PartRem[33][7] ), .B(
        net32242), .CI(\u_div/CryTmp[32][7] ), .CO(\u_div/CryTmp[32][8] ), .S(
        \u_div/SumTmp[32][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_8  ( .A(\u_div/PartRem[33][8] ), .B(
        net32200), .CI(n254), .CO(\u_div/CryTmp[32][9] ), .S(
        \u_div/SumTmp[32][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_9  ( .A(\u_div/PartRem[33][9] ), .B(
        net32186), .CI(\u_div/CryTmp[32][9] ), .CO(\u_div/CryTmp[32][10] ), 
        .S(\u_div/SumTmp[32][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_10  ( .A(\u_div/PartRem[33][10] ), .B(
        net32140), .CI(\u_div/CryTmp[32][10] ), .CO(\u_div/CryTmp[32][11] ), 
        .S(\u_div/SumTmp[32][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_11  ( .A(n326), .B(n445), .CI(net49055), 
        .CO(\u_div/CryTmp[32][12] ), .S(\u_div/SumTmp[32][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_12  ( .A(\u_div/PartRem[33][12] ), .B(
        net32088), .CI(\u_div/CryTmp[32][12] ), .CO(\u_div/CryTmp[32][13] ), 
        .S(\u_div/SumTmp[32][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_32_13  ( .A(\u_div/PartRem[33][13] ), .B(
        net32078), .CI(n230), .CO(\u_div/CryTmp[32][14] ), .S(
        \u_div/SumTmp[32][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_2  ( .A(\u_div/PartRem[32][2] ), .B(
        net32366), .CI(\u_div/CryTmp[31][2] ), .CO(\u_div/CryTmp[31][3] ), .S(
        \u_div/SumTmp[31][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_3  ( .A(\u_div/PartRem[32][3] ), .B(
        net32338), .CI(\u_div/CryTmp[31][3] ), .CO(\u_div/CryTmp[31][4] ), .S(
        \u_div/SumTmp[31][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_4  ( .A(\u_div/PartRem[32][4] ), .B(
        net32314), .CI(\u_div/CryTmp[31][4] ), .CO(\u_div/CryTmp[31][5] ), .S(
        \u_div/SumTmp[31][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_6  ( .A(\u_div/PartRem[32][6] ), .B(
        net32254), .CI(\u_div/CryTmp[31][6] ), .CO(\u_div/CryTmp[31][7] ), .S(
        \u_div/SumTmp[31][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_7  ( .A(\u_div/PartRem[32][7] ), .B(
        net32226), .CI(\u_div/CryTmp[31][7] ), .CO(\u_div/CryTmp[31][8] ), .S(
        \u_div/SumTmp[31][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_8  ( .A(\u_div/PartRem[32][8] ), .B(
        net32200), .CI(n437), .CO(\u_div/CryTmp[31][9] ), .S(
        \u_div/SumTmp[31][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_9  ( .A(\u_div/PartRem[32][9] ), .B(
        net32186), .CI(\u_div/CryTmp[31][9] ), .CO(\u_div/CryTmp[31][10] ), 
        .S(\u_div/SumTmp[31][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_10  ( .A(\u_div/PartRem[32][10] ), .B(
        \u_div/CryTmp[31][10] ), .CI(net32140), .CO(\u_div/CryTmp[31][11] ), 
        .S(\u_div/SumTmp[31][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_12  ( .A(\u_div/PartRem[32][12] ), .B(
        net32088), .CI(n439), .CO(\u_div/CryTmp[31][13] ), .S(
        \u_div/SumTmp[31][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_13  ( .A(\u_div/PartRem[32][13] ), .B(
        net32078), .CI(n61), .CO(\u_div/CryTmp[31][14] ), .S(
        \u_div/SumTmp[31][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_14  ( .A(\u_div/PartRem[32][14] ), .B(
        net32046), .CI(\u_div/CryTmp[31][14] ), .CO(\u_div/CryTmp[31][15] ), 
        .S(\u_div/SumTmp[31][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_1  ( .A(\u_div/PartRem[31][1] ), .B(
        net32386), .CI(\u_div/CryTmp[30][1] ), .CO(\u_div/CryTmp[30][2] ), .S(
        \u_div/SumTmp[30][1] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_30_2  ( .A(\u_div/PartRem[31][2] ), .B(
        net32366), .CI(\u_div/CryTmp[30][2] ), .CO(\u_div/CryTmp[30][3] ), .S(
        \u_div/SumTmp[30][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_3  ( .A(\u_div/PartRem[31][3] ), .B(
        net32338), .CI(n454), .CO(\u_div/CryTmp[30][4] ), .S(
        \u_div/SumTmp[30][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_4  ( .A(\u_div/PartRem[31][4] ), .B(
        net32314), .CI(\u_div/CryTmp[30][4] ), .CO(\u_div/CryTmp[30][5] ), .S(
        \u_div/SumTmp[30][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_5  ( .A(\u_div/PartRem[31][5] ), .B(
        net32284), .CI(n456), .CO(\u_div/CryTmp[30][6] ), .S(
        \u_div/SumTmp[30][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_6  ( .A(\u_div/PartRem[31][6] ), .B(
        net32254), .CI(\u_div/CryTmp[30][6] ), .CO(\u_div/CryTmp[30][7] ), .S(
        \u_div/SumTmp[30][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_7  ( .A(\u_div/PartRem[31][7] ), .B(
        net32222), .CI(\u_div/CryTmp[30][7] ), .CO(\u_div/CryTmp[30][8] ), .S(
        \u_div/SumTmp[30][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_8  ( .A(\u_div/PartRem[31][8] ), .B(
        net32200), .CI(\u_div/CryTmp[30][8] ), .CO(\u_div/CryTmp[30][9] ), .S(
        \u_div/SumTmp[30][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_9  ( .A(\u_div/PartRem[31][9] ), .B(
        net32166), .CI(\u_div/CryTmp[30][9] ), .CO(\u_div/CryTmp[30][10] ), 
        .S(\u_div/SumTmp[30][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_10  ( .A(\u_div/PartRem[31][10] ), .B(
        net32140), .CI(\u_div/CryTmp[30][10] ), .CO(\u_div/CryTmp[30][11] ), 
        .S(\u_div/SumTmp[30][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_11  ( .A(\u_div/PartRem[31][11] ), .B(
        net49055), .CI(\u_div/CryTmp[30][11] ), .CO(\u_div/CryTmp[30][12] ), 
        .S(\u_div/SumTmp[30][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_12  ( .A(\u_div/PartRem[31][12] ), .B(
        net32088), .CI(\u_div/CryTmp[30][12] ), .CO(\u_div/CryTmp[30][13] ), 
        .S(\u_div/SumTmp[30][12] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_13  ( .A(n452), .B(net32078), .CI(n443), 
        .CO(\u_div/CryTmp[30][14] ), .S(\u_div/SumTmp[30][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_14  ( .A(\u_div/PartRem[31][14] ), .B(
        net32046), .CI(\u_div/CryTmp[30][14] ), .CO(\u_div/CryTmp[30][15] ), 
        .S(\u_div/SumTmp[30][14] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_15  ( .A(\u_div/PartRem[31][15] ), .B(
        net32016), .CI(\u_div/CryTmp[30][15] ), .CO(\u_div/CryTmp[30][16] ), 
        .S(\u_div/SumTmp[30][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_30_16  ( .A(n448), .B(net31982), .CI(
        \u_div/PartRem[31][16] ), .CO(\u_div/CryTmp[30][17] ), .S(
        \u_div/SumTmp[30][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_44_1  ( .A(\u_div/CryTmp[44][1] ), .B(
        net32382), .CI(\u_div/PartRem[45][1] ), .CO(\u_div/CryTmp[44][2] ), 
        .S(\u_div/SumTmp[44][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_44_2  ( .A(\u_div/PartRem[45][2] ), .B(
        net32368), .CI(\u_div/CryTmp[44][2] ), .CO(\u_div/CryTmp[44][3] ), .S(
        \u_div/SumTmp[44][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_43_1  ( .A(\u_div/PartRem[44][1] ), .B(
        net32382), .CI(\u_div/CryTmp[43][1] ), .CO(\u_div/CryTmp[43][2] ), .S(
        \u_div/SumTmp[43][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_43_2  ( .A(\u_div/PartRem[44][2] ), .B(
        net32368), .CI(n308), .CO(\u_div/CryTmp[43][3] ), .S(
        \u_div/SumTmp[43][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_43_3  ( .A(\u_div/PartRem[44][3] ), .B(
        net32354), .CI(\u_div/CryTmp[43][3] ), .CO(\u_div/CryTmp[43][4] ), .S(
        \u_div/SumTmp[43][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_42_1  ( .A(net32382), .B(
        \u_div/PartRem[43][1] ), .CI(\u_div/CryTmp[42][1] ), .CO(
        \u_div/CryTmp[42][2] ), .S(\u_div/SumTmp[42][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_42_2  ( .A(\u_div/PartRem[43][2] ), .B(
        net32368), .CI(\u_div/CryTmp[42][2] ), .CO(\u_div/CryTmp[42][3] ), .S(
        \u_div/SumTmp[42][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_42_3  ( .A(\u_div/PartRem[43][3] ), .B(
        net32354), .CI(\u_div/CryTmp[42][3] ), .CO(\u_div/CryTmp[42][4] ), .S(
        \u_div/SumTmp[42][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_42_4  ( .A(\u_div/PartRem[43][4] ), .B(
        net32326), .CI(\u_div/CryTmp[42][4] ), .CO(\u_div/CryTmp[42][5] ), .S(
        \u_div/SumTmp[42][4] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_41_1  ( .A(n377), .B(net32382), .CI(
        \u_div/CryTmp[41][1] ), .CO(\u_div/CryTmp[41][2] ), .S(
        \u_div/SumTmp[41][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_41_2  ( .A(n168), .B(net32368), .CI(n384), 
        .CO(\u_div/CryTmp[41][3] ), .S(\u_div/SumTmp[41][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_41_3  ( .A(\u_div/PartRem[42][3] ), .B(
        net32354), .CI(\u_div/CryTmp[41][3] ), .CO(\u_div/CryTmp[41][4] ), .S(
        \u_div/SumTmp[41][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_41_4  ( .A(\u_div/PartRem[42][4] ), .B(
        net32326), .CI(n218), .CO(\u_div/CryTmp[41][5] ), .S(
        \u_div/SumTmp[41][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_41_5  ( .A(\u_div/PartRem[42][5] ), .B(
        net32302), .CI(\u_div/CryTmp[41][5] ), .CO(\u_div/CryTmp[41][6] ), .S(
        \u_div/SumTmp[41][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_40_1  ( .A(\u_div/PartRem[41][1] ), .B(
        net32382), .CI(\u_div/CryTmp[40][1] ), .CO(\u_div/CryTmp[40][2] ), .S(
        \u_div/SumTmp[40][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_40_2  ( .A(\u_div/PartRem[41][2] ), .B(
        net32368), .CI(\u_div/CryTmp[40][2] ), .CO(\u_div/CryTmp[40][3] ), .S(
        \u_div/SumTmp[40][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_40_3  ( .A(\u_div/PartRem[41][3] ), .B(
        net32354), .CI(\u_div/CryTmp[40][3] ), .CO(\u_div/CryTmp[40][4] ), .S(
        \u_div/SumTmp[40][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_40_4  ( .A(\u_div/PartRem[41][4] ), .B(
        net32326), .CI(\u_div/CryTmp[40][4] ), .CO(\u_div/CryTmp[40][5] ), .S(
        \u_div/SumTmp[40][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_40_5  ( .A(\u_div/PartRem[41][5] ), .B(
        net32302), .CI(\u_div/CryTmp[40][5] ), .CO(\u_div/CryTmp[40][6] ), .S(
        \u_div/SumTmp[40][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_40_6  ( .A(\u_div/PartRem[41][6] ), .B(
        net32272), .CI(\u_div/CryTmp[40][6] ), .CO(\u_div/CryTmp[40][7] ), .S(
        \u_div/SumTmp[40][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_39_7  ( .A(\u_div/PartRem[40][7] ), .B(
        net32242), .CI(\u_div/CryTmp[39][7] ), .CO(\u_div/CryTmp[39][8] ), .S(
        \u_div/SumTmp[39][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_39_1  ( .A(\u_div/PartRem[40][1] ), .B(
        net32382), .CI(\u_div/CryTmp[39][1] ), .CO(\u_div/CryTmp[39][2] ), .S(
        \u_div/SumTmp[39][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_39_2  ( .A(\u_div/PartRem[40][2] ), .B(
        net32368), .CI(n380), .CO(\u_div/CryTmp[39][3] ), .S(
        \u_div/SumTmp[39][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_39_3  ( .A(\u_div/PartRem[40][3] ), .B(
        net32354), .CI(\u_div/CryTmp[39][3] ), .CO(\u_div/CryTmp[39][4] ), .S(
        \u_div/SumTmp[39][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_39_4  ( .A(\u_div/PartRem[40][4] ), .B(
        net32326), .CI(\u_div/CryTmp[39][4] ), .CO(\u_div/CryTmp[39][5] ), .S(
        \u_div/SumTmp[39][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_39_5  ( .A(\u_div/PartRem[40][5] ), .B(
        net32302), .CI(\u_div/CryTmp[39][5] ), .CO(\u_div/CryTmp[39][6] ), .S(
        \u_div/SumTmp[39][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_39_6  ( .A(\u_div/PartRem[40][6] ), .B(
        net32272), .CI(\u_div/CryTmp[39][6] ), .CO(\u_div/CryTmp[39][7] ), .S(
        \u_div/SumTmp[39][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_1  ( .A(\u_div/PartRem[39][1] ), .B(
        net32382), .CI(\u_div/CryTmp[38][1] ), .CO(\u_div/CryTmp[38][2] ), .S(
        \u_div/SumTmp[38][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_2  ( .A(\u_div/PartRem[39][2] ), .B(
        net32368), .CI(\u_div/CryTmp[38][2] ), .CO(\u_div/CryTmp[38][3] ), .S(
        \u_div/SumTmp[38][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_3  ( .A(\u_div/PartRem[39][3] ), .B(
        net32354), .CI(\u_div/CryTmp[38][3] ), .CO(\u_div/CryTmp[38][4] ), .S(
        \u_div/SumTmp[38][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_4  ( .A(\u_div/PartRem[39][4] ), .B(
        net32326), .CI(n65), .CO(\u_div/CryTmp[38][5] ), .S(
        \u_div/SumTmp[38][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_5  ( .A(\u_div/PartRem[39][5] ), .B(
        net32302), .CI(\u_div/CryTmp[38][5] ), .CO(\u_div/CryTmp[38][6] ), .S(
        \u_div/SumTmp[38][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_6  ( .A(\u_div/PartRem[39][6] ), .B(
        net32272), .CI(\u_div/CryTmp[38][6] ), .CO(\u_div/CryTmp[38][7] ), .S(
        \u_div/SumTmp[38][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_7  ( .A(\u_div/PartRem[39][7] ), .B(
        net32242), .CI(n382), .CO(\u_div/CryTmp[38][8] ), .S(
        \u_div/SumTmp[38][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_38_8  ( .A(\u_div/PartRem[39][8] ), .B(
        net32212), .CI(\u_div/CryTmp[38][8] ), .CO(\u_div/CryTmp[38][9] ), .S(
        \u_div/SumTmp[38][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_1  ( .A(\u_div/PartRem[38][1] ), .B(
        net32382), .CI(\u_div/CryTmp[37][1] ), .CO(\u_div/CryTmp[37][2] ), .S(
        \u_div/SumTmp[37][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_37_2  ( .A(net46015), .B(net32368), .CI(
        \u_div/CryTmp[37][2] ), .CO(\u_div/CryTmp[37][3] ), .S(
        \u_div/SumTmp[37][2] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_17  ( .A(\u_div/PartRem[2][17] ), .B(
        net31964), .CI(\u_div/CryTmp[1][17] ), .CO(\u_div/CryTmp[1][18] ), .S(
        \u_div/SumTmp[1][17] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_21_13  ( .A(\u_div/PartRem[22][13] ), .B(
        net32066), .CI(\u_div/CryTmp[21][13] ), .CO(\u_div/CryTmp[21][14] ), 
        .S(\u_div/SumTmp[21][13] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_25_18  ( .A(\u_div/PartRem[26][18] ), .B(
        net31938), .CI(n517), .CO(\u_div/CryTmp[25][19] ), .S(
        \u_div/SumTmp[25][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_20  ( .A(\u_div/PartRem[24][20] ), .B(
        net31884), .CI(\u_div/CryTmp[23][20] ), .CO(\u_div/CryTmp[23][21] ), 
        .S(\u_div/SumTmp[23][20] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_17_6  ( .A(\u_div/PartRem[18][6] ), .B(
        net32252), .CI(\u_div/CryTmp[17][6] ), .CO(\u_div/CryTmp[17][7] ), .S(
        \u_div/SumTmp[17][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_11  ( .A(\u_div/PartRem[36][11] ), .B(
        net49055), .CI(n961), .CO(\u_div/CryTmp[35][12] ), .S(
        \u_div/SumTmp[35][11] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_36_9  ( .A(\u_div/PartRem[37][9] ), .B(
        net32186), .CI(n284), .CO(\u_div/CryTmp[36][10] ), .S(
        \u_div/SumTmp[36][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_25_21  ( .A(\u_div/PartRem[26][21] ), .B(
        net31856), .CI(n294), .CO(\u_div/CryTmp[25][22] ), .S(
        \u_div/SumTmp[25][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_22  ( .A(\u_div/PartRem[2][22] ), .B(
        net31826), .CI(n226), .CO(\u_div/CryTmp[1][23] ), .S(
        \u_div/SumTmp[1][22] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_20  ( .A(\u_div/PartRem[1][20] ), .B(
        net31882), .CI(\u_div/CryTmp[0][20] ), .CO(\u_div/CryTmp[0][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_21  ( .A(\u_div/PartRem[4][21] ), .B(
        net31854), .CI(\u_div/CryTmp[3][21] ), .CO(\u_div/CryTmp[3][22] ), .S(
        \u_div/SumTmp[3][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_21  ( .A(\u_div/PartRem[10][21] ), .B(
        net31854), .CI(\u_div/CryTmp[9][21] ), .CO(\u_div/CryTmp[9][22] ), .S(
        \u_div/SumTmp[9][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_21  ( .A(\u_div/PartRem[13][21] ), .B(
        net31856), .CI(\u_div/CryTmp[12][21] ), .CO(\u_div/CryTmp[12][22] ), 
        .S(\u_div/SumTmp[12][21] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_0_18  ( .A(\u_div/PartRem[1][18] ), .B(
        net31940), .CI(n946), .CO(\u_div/CryTmp[0][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_36_6  ( .A(\u_div/PartRem[37][6] ), .B(
        net32272), .CI(\u_div/CryTmp[36][6] ), .CO(\u_div/CryTmp[36][7] ), .S(
        \u_div/SumTmp[36][6] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_8  ( .A(\u_div/PartRem[35][8] ), .B(
        net32200), .CI(\u_div/CryTmp[34][8] ), .CO(\u_div/CryTmp[34][9] ), .S(
        \u_div/SumTmp[34][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_19  ( .A(n857), .B(net31910), .CI(
        \u_div/CryTmp[3][19] ), .CO(\u_div/CryTmp[3][20] ), .S(
        \u_div/SumTmp[3][19] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_11_18  ( .A(\u_div/PartRem[12][18] ), .B(
        net31940), .CI(\u_div/CryTmp[11][18] ), .CO(\u_div/CryTmp[11][19] ), 
        .S(\u_div/SumTmp[11][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_6_17  ( .A(\u_div/PartRem[7][17] ), .B(
        net31962), .CI(\u_div/CryTmp[6][17] ), .CO(\u_div/CryTmp[6][18] ), .S(
        \u_div/SumTmp[6][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_13  ( .A(\u_div/PartRem[2][13] ), .B(
        net32068), .CI(n914), .CO(\u_div/CryTmp[1][14] ), .S(
        \u_div/SumTmp[1][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_10_16  ( .A(\u_div/PartRem[11][16] ), .B(
        net31984), .CI(n304), .CO(\u_div/CryTmp[10][17] ), .S(
        \u_div/SumTmp[10][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_23_16  ( .A(\u_div/PartRem[24][16] ), .B(
        net31982), .CI(n73), .CO(\u_div/CryTmp[23][17] ), .S(
        \u_div/SumTmp[23][16] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_15  ( .A(\u_div/PartRem[13][15] ), .B(
        net32014), .CI(\u_div/CryTmp[12][15] ), .CO(\u_div/CryTmp[12][16] ), 
        .S(\u_div/SumTmp[12][15] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_1_8  ( .A(n951), .B(net32196), .CI(n999), 
        .CO(\u_div/CryTmp[1][9] ), .S(\u_div/SumTmp[1][8] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_3_11  ( .A(\u_div/PartRem[4][11] ), .B(
        net32118), .CI(\u_div/CryTmp[3][11] ), .CO(\u_div/CryTmp[3][12] ), .S(
        \u_div/SumTmp[3][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_8_13  ( .A(\u_div/PartRem[9][13] ), .B(
        net32068), .CI(\u_div/CryTmp[8][13] ), .CO(\u_div/CryTmp[8][14] ), .S(
        \u_div/SumTmp[8][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_5  ( .A(\u_div/PartRem[32][5] ), .B(
        net32284), .CI(\u_div/CryTmp[31][5] ), .CO(\u_div/CryTmp[31][6] ), .S(
        \u_div/SumTmp[31][5] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_15_11  ( .A(\u_div/PartRem[16][11] ), .B(
        net32116), .CI(\u_div/CryTmp[15][11] ), .CO(\u_div/CryTmp[15][12] ), 
        .S(\u_div/SumTmp[15][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_4_4  ( .A(\u_div/PartRem[5][4] ), .B(
        net32310), .CI(\u_div/CryTmp[4][4] ), .CO(\u_div/CryTmp[4][5] ), .S(
        \u_div/SumTmp[4][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_7  ( .A(\u_div/PartRem[27][7] ), .B(
        net32222), .CI(\u_div/CryTmp[26][7] ), .CO(\u_div/CryTmp[26][8] ), .S(
        \u_div/SumTmp[26][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_9_4  ( .A(\u_div/PartRem[10][4] ), .B(
        net32310), .CI(\u_div/CryTmp[9][4] ), .CO(\u_div/CryTmp[9][5] ), .S(
        \u_div/SumTmp[9][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_21_4  ( .A(\u_div/PartRem[22][4] ), .B(
        net32312), .CI(\u_div/CryTmp[21][4] ), .CO(\u_div/CryTmp[21][5] ), .S(
        \u_div/SumTmp[21][4] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_34_10  ( .A(\u_div/PartRem[35][10] ), .B(
        net32140), .CI(\u_div/CryTmp[34][10] ), .CO(\u_div/CryTmp[34][11] ), 
        .S(\u_div/SumTmp[34][10] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_12_20  ( .A(\u_div/PartRem[13][20] ), .B(
        net31884), .CI(\u_div/CryTmp[12][20] ), .CO(\u_div/CryTmp[12][21] ), 
        .S(\u_div/SumTmp[12][20] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_18  ( .A(\u_div/PartRem[18][18] ), .B(
        net31938), .CI(\u_div/CryTmp[17][18] ), .CO(\u_div/CryTmp[17][19] ), 
        .S(\u_div/SumTmp[17][18] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_13_17  ( .A(\u_div/PartRem[14][17] ), .B(
        net31962), .CI(\u_div/CryTmp[13][17] ), .CO(\u_div/CryTmp[13][18] ), 
        .S(\u_div/SumTmp[13][17] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_13  ( .A(\u_div/PartRem[20][13] ), .B(
        net32066), .CI(\u_div/CryTmp[19][13] ), .CO(\u_div/CryTmp[19][14] ), 
        .S(\u_div/SumTmp[19][13] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_19_9  ( .A(\u_div/PartRem[20][9] ), .B(
        net32166), .CI(\u_div/CryTmp[19][9] ), .CO(\u_div/CryTmp[19][10] ), 
        .S(\u_div/SumTmp[19][9] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_17_7  ( .A(\u_div/PartRem[18][7] ), .B(
        net32222), .CI(n628), .CO(\u_div/CryTmp[17][8] ), .S(
        \u_div/SumTmp[17][7] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_26_3  ( .A(\u_div/PartRem[27][3] ), .B(
        net32338), .CI(\u_div/CryTmp[26][3] ), .CO(\u_div/CryTmp[26][4] ), .S(
        \u_div/SumTmp[26][3] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_24_1  ( .A(net41045), .B(net32386), .CI(
        \u_div/CryTmp[24][1] ), .CO(\u_div/CryTmp[24][2] ), .S(
        \u_div/SumTmp[24][1] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_31_11  ( .A(\u_div/PartRem[32][11] ), .B(
        net49055), .CI(\u_div/CryTmp[31][11] ), .CO(\u_div/CryTmp[31][12] ), 
        .S(\u_div/SumTmp[31][11] ) );
  FADDX1_RVT \u_div/u_fa_PartRem_0_35_5  ( .A(\u_div/PartRem[36][5] ), .B(
        net32284), .CI(\u_div/CryTmp[35][5] ), .CO(\u_div/CryTmp[35][6] ), .S(
        \u_div/SumTmp[35][5] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_4_18  ( .A(\u_div/PartRem[5][18] ), .B(
        net31940), .CI(\u_div/CryTmp[4][18] ), .CO(\u_div/CryTmp[4][19] ), .S(
        \u_div/SumTmp[4][18] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_26_9  ( .A(\u_div/PartRem[27][9] ), .B(
        net32168), .CI(\u_div/CryTmp[26][9] ), .CO(\u_div/CryTmp[26][10] ), 
        .S(\u_div/SumTmp[26][9] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_29_9  ( .A(\u_div/PartRem[30][9] ), .B(
        net32166), .CI(\u_div/CryTmp[29][9] ), .CO(\u_div/CryTmp[29][10] ), 
        .S(\u_div/SumTmp[29][9] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_1_21  ( .A(\u_div/PartRem[2][21] ), .B(
        net31854), .CI(\u_div/CryTmp[1][21] ), .CO(\u_div/CryTmp[1][22] ), .S(
        \u_div/SumTmp[1][21] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_25_10  ( .A(\u_div/PartRem[26][10] ), .B(
        net32140), .CI(\u_div/CryTmp[25][10] ), .CO(\u_div/CryTmp[25][11] ), 
        .S(\u_div/SumTmp[25][10] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_5_21  ( .A(\u_div/PartRem[6][21] ), .B(
        net31854), .CI(\u_div/CryTmp[5][21] ), .CO(\u_div/CryTmp[5][22] ), .S(
        \u_div/SumTmp[5][21] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_22_14  ( .A(\u_div/PartRem[23][14] ), .B(
        net32044), .CI(\u_div/CryTmp[22][14] ), .CO(\u_div/CryTmp[22][15] ), 
        .S(\u_div/SumTmp[22][14] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_3_5  ( .A(\u_div/PartRem[4][5] ), .B(
        net32280), .CI(\u_div/CryTmp[3][5] ), .CO(\u_div/CryTmp[3][6] ), .S(
        \u_div/SumTmp[3][5] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_12_18  ( .A(\u_div/PartRem[13][18] ), .B(
        net31940), .CI(\u_div/CryTmp[12][18] ), .CO(\u_div/CryTmp[12][19] ), 
        .S(\u_div/SumTmp[12][18] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_21_6  ( .A(\u_div/PartRem[22][6] ), .B(
        net32252), .CI(\u_div/CryTmp[21][6] ), .CO(\u_div/CryTmp[21][7] ), .S(
        \u_div/SumTmp[21][6] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_9_13  ( .A(\u_div/PartRem[10][13] ), .B(
        net32068), .CI(\u_div/CryTmp[9][13] ), .CO(\u_div/CryTmp[9][14] ), .S(
        \u_div/SumTmp[9][13] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_35_10  ( .A(\u_div/CryTmp[35][10] ), .B(
        net32140), .CI(\u_div/PartRem[36][10] ), .CO(\u_div/CryTmp[35][11] ), 
        .S(\u_div/SumTmp[35][10] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_20_14  ( .A(net32044), .B(
        \u_div/PartRem[21][14] ), .CI(\u_div/CryTmp[20][14] ), .CO(
        \u_div/CryTmp[20][15] ), .S(\u_div/SumTmp[20][14] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_17_21  ( .A(\u_div/PartRem[18][21] ), .B(
        \u_div/CryTmp[17][21] ), .CI(net31856), .CO(\u_div/CryTmp[17][22] ), 
        .S(\u_div/SumTmp[17][21] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_14_15  ( .A(\u_div/PartRem[15][15] ), .B(
        net32014), .CI(\u_div/CryTmp[14][15] ), .CO(\u_div/CryTmp[14][16] ), 
        .S(\u_div/SumTmp[14][15] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_16_4  ( .A(\u_div/PartRem[17][4] ), .B(
        \u_div/CryTmp[16][4] ), .CI(net32312), .CO(\u_div/CryTmp[16][5] ), .S(
        \u_div/SumTmp[16][4] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_28_16  ( .A(\u_div/PartRem[29][16] ), .B(
        net31982), .CI(n934), .CO(\u_div/CryTmp[28][17] ), .S(
        \u_div/SumTmp[28][16] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_10_19  ( .A(\u_div/PartRem[11][19] ), .B(
        net31910), .CI(\u_div/CryTmp[10][19] ), .CO(\u_div/CryTmp[10][20] ), 
        .S(\u_div/SumTmp[10][19] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_15_19  ( .A(\u_div/PartRem[16][19] ), .B(
        net31912), .CI(\u_div/CryTmp[15][19] ), .CO(\u_div/CryTmp[15][20] ), 
        .S(\u_div/SumTmp[15][19] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_3_12  ( .A(\u_div/PartRem[4][12] ), .B(n863), .CI(net32092), .CO(\u_div/CryTmp[3][13] ), .S(\u_div/SumTmp[3][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_23_21  ( .A(\u_div/PartRem[24][21] ), .B(
        net31856), .CI(\u_div/CryTmp[23][21] ), .CO(\u_div/CryTmp[23][22] ), 
        .S(\u_div/SumTmp[23][21] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_18_22  ( .A(\u_div/PartRem[19][22] ), .B(
        net31828), .CI(\u_div/CryTmp[18][22] ), .CO(\u_div/CryTmp[18][23] ), 
        .S(\u_div/SumTmp[18][22] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_13_22  ( .A(\u_div/PartRem[14][22] ), .B(
        net31828), .CI(\u_div/CryTmp[13][22] ), .CO(\u_div/CryTmp[13][23] ), 
        .S(\u_div/SumTmp[13][22] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_33_12  ( .A(\u_div/PartRem[34][12] ), .B(
        net32088), .CI(\u_div/CryTmp[33][12] ), .CO(\u_div/CryTmp[33][13] ), 
        .S(\u_div/SumTmp[33][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_11_9  ( .A(\u_div/PartRem[12][9] ), .B(
        net32168), .CI(\u_div/CryTmp[11][9] ), .CO(\u_div/CryTmp[11][10] ), 
        .S(\u_div/SumTmp[11][9] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_45_1  ( .A(\u_div/CryTmp[45][1] ), .B(
        net32384), .CI(\u_div/PartRem[46][1] ), .CO(\u_div/CryTmp[45][2] ), 
        .S(\u_div/SumTmp[45][1] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_31_1  ( .A(\u_div/PartRem[32][1] ), .B(
        net32386), .CI(\u_div/CryTmp[31][1] ), .CO(\u_div/CryTmp[31][2] ), .S(
        \u_div/SumTmp[31][1] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_20_12  ( .A(n123), .B(net32090), .CI(n160), 
        .CO(\u_div/CryTmp[20][13] ), .S(\u_div/SumTmp[20][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_34_12  ( .A(\u_div/PartRem[35][12] ), .B(
        net32088), .CI(\u_div/CryTmp[34][12] ), .CO(\u_div/CryTmp[34][13] ), 
        .S(\u_div/SumTmp[34][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_4_11  ( .A(\u_div/PartRem[5][11] ), .B(
        net32118), .CI(\u_div/CryTmp[4][11] ), .CO(\u_div/CryTmp[4][12] ), .S(
        \u_div/SumTmp[4][11] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_28_12  ( .A(\u_div/PartRem[29][12] ), .B(
        net32088), .CI(\u_div/CryTmp[28][12] ), .CO(\u_div/CryTmp[28][13] ), 
        .S(\u_div/SumTmp[28][12] ) );
  FADDX2_RVT \u_div/u_fa_PartRem_0_27_8  ( .A(\u_div/PartRem[28][8] ), .B(
        net32200), .CI(\u_div/CryTmp[27][8] ), .CO(\u_div/CryTmp[27][9] ), .S(
        \u_div/SumTmp[27][8] ) );
  INVX1_RVT U1 ( .A(net38350), .Y(net50726) );
  INVX4_RVT U2 ( .A(net50727), .Y(net42040) );
  IBUFFX4_RVT U3 ( .A(net40598), .Y(net38350) );
  IBUFFX16_RVT U4 ( .A(\u_div/CryTmp[8][8] ), .Y(n1) );
  INVX2_RVT U5 ( .A(n1), .Y(n2) );
  INVX0_RVT U6 ( .A(net29664), .Y(\u_div/PartRem[7][16] ) );
  NOR2X4_RVT U7 ( .A1(\u_div/CryTmp[21][24] ), .A2(\u_div/PartRem[22][24] ), 
        .Y(net38342) );
  INVX1_RVT U8 ( .A(net45183), .Y(net45594) );
  IBUFFX4_RVT U9 ( .A(net45183), .Y(net45597) );
  INVX8_RVT U10 ( .A(net45183), .Y(n842) );
  INVX1_RVT U11 ( .A(\u_div/CryTmp[14][21] ), .Y(net48638) );
  IBUFFX16_RVT U12 ( .A(\u_div/SumTmp[15][17] ), .Y(net30977) );
  IBUFFX4_RVT U13 ( .A(net38341), .Y(n3) );
  NBUFFX8_RVT U14 ( .A(net38341), .Y(n4) );
  INVX8_RVT U15 ( .A(n4), .Y(n5) );
  IBUFFX4_RVT U16 ( .A(n4), .Y(n6) );
  IBUFFX4_RVT U17 ( .A(n4), .Y(n7) );
  INVX1_RVT U18 ( .A(n3), .Y(n8) );
  INVX1_RVT U19 ( .A(n3), .Y(n9) );
  INVX1_RVT U20 ( .A(n3), .Y(n10) );
  INVX0_RVT U21 ( .A(n8), .Y(n11) );
  INVX0_RVT U22 ( .A(n8), .Y(n12) );
  INVX0_RVT U23 ( .A(n8), .Y(n13) );
  INVX0_RVT U24 ( .A(n8), .Y(n14) );
  INVX0_RVT U25 ( .A(n9), .Y(n15) );
  INVX0_RVT U26 ( .A(n9), .Y(n16) );
  INVX0_RVT U27 ( .A(n9), .Y(n17) );
  INVX0_RVT U28 ( .A(n9), .Y(n18) );
  INVX1_RVT U29 ( .A(n10), .Y(n19) );
  INVX0_RVT U30 ( .A(n10), .Y(n20) );
  INVX0_RVT U31 ( .A(n10), .Y(quotient[16]) );
  INVX1_RVT U32 ( .A(n10), .Y(n22) );
  NOR2X1_RVT U33 ( .A1(\u_div/PartRem[17][24] ), .A2(\u_div/CryTmp[16][24] ), 
        .Y(net38341) );
  IBUFFX4_RVT U34 ( .A(n729), .Y(\u_div/PartRem[12][10] ) );
  IBUFFX16_RVT U35 ( .A(\u_div/CryTmp[15][3] ), .Y(n23) );
  INVX4_RVT U36 ( .A(n23), .Y(n24) );
  INVX2_RVT U37 ( .A(n1142), .Y(\u_div/PartRem[2][23] ) );
  IBUFFX4_RVT U38 ( .A(net30658), .Y(\u_div/PartRem[16][18] ) );
  INVX4_RVT U39 ( .A(n291), .Y(n25) );
  IBUFFX4_RVT U40 ( .A(n25), .Y(n26) );
  IBUFFX2_RVT U41 ( .A(\u_div/PartRem[27][13] ), .Y(n27) );
  IBUFFX4_RVT U42 ( .A(n27), .Y(n28) );
  IBUFFX16_RVT U43 ( .A(net30000), .Y(\u_div/PartRem[27][13] ) );
  MUX21X2_RVT U44 ( .A1(n798), .A2(n830), .S0(net44755), .Y(n816) );
  IBUFFX32_RVT U45 ( .A(\u_div/SumTmp[5][14] ), .Y(n830) );
  MUX21X2_RVT U46 ( .A1(net29667), .A2(net30384), .S0(net45257), .Y(n798) );
  IBUFFX4_RVT U47 ( .A(net30853), .Y(net45940) );
  NBUFFX2_RVT U48 ( .A(net30501), .Y(n29) );
  INVX1_RVT U49 ( .A(\u_div/SumTmp[33][9] ), .Y(net30501) );
  IBUFFX4_RVT U50 ( .A(\u_div/PartRem[14][10] ), .Y(n30) );
  INVX4_RVT U51 ( .A(n30), .Y(n31) );
  INVX4_RVT U52 ( .A(\u_div/PartRem[23][16] ), .Y(n32) );
  INVX1_RVT U53 ( .A(n32), .Y(n33) );
  IBUFFX4_RVT U54 ( .A(n550), .Y(\u_div/PartRem[21][15] ) );
  NBUFFX8_RVT U55 ( .A(net31184), .Y(n34) );
  IBUFFX4_RVT U56 ( .A(\u_div/CryTmp[11][17] ), .Y(n35) );
  INVX2_RVT U57 ( .A(n35), .Y(n36) );
  IBUFFX16_RVT U58 ( .A(\u_div/SumTmp[13][8] ), .Y(net31184) );
  MUX21X2_RVT U59 ( .A1(n1023), .A2(n1152), .S0(net32520), .Y(net29665) );
  INVX32_RVT U60 ( .A(n1023), .Y(\u_div/PartRem[8][14] ) );
  MUX21X2_RVT U61 ( .A1(net29616), .A2(net30366), .S0(net40719), .Y(n1023) );
  MUX21X2_RVT U62 ( .A1(n1024), .A2(n1155), .S0(net46859), .Y(net29666) );
  INVX32_RVT U63 ( .A(n1024), .Y(\u_div/PartRem[8][13] ) );
  MUX21X2_RVT U64 ( .A1(net29617), .A2(net30376), .S0(net40719), .Y(n1024) );
  MUX21X2_RVT U65 ( .A1(n1025), .A2(n1158), .S0(net46859), .Y(net29667) );
  INVX32_RVT U66 ( .A(n1025), .Y(\u_div/PartRem[8][12] ) );
  MUX21X2_RVT U67 ( .A1(net29618), .A2(net30386), .S0(net40719), .Y(n1025) );
  IBUFFX4_RVT U68 ( .A(\u_div/PartRem[7][12] ), .Y(n37) );
  INVX1_RVT U69 ( .A(n37), .Y(n38) );
  IBUFFX4_RVT U70 ( .A(net29668), .Y(\u_div/PartRem[7][12] ) );
  IBUFFX4_RVT U71 ( .A(\u_div/PartRem[34][13] ), .Y(n39) );
  INVX1_RVT U72 ( .A(n39), .Y(n40) );
  IBUFFX16_RVT U73 ( .A(net29872), .Y(\u_div/PartRem[34][13] ) );
  IBUFFX4_RVT U74 ( .A(\u_div/SumTmp[28][12] ), .Y(n1183) );
  MUX21X1_RVT U75 ( .A1(net29668), .A2(net30394), .S0(net45257), .Y(n799) );
  IBUFFX4_RVT U76 ( .A(n591), .Y(\u_div/PartRem[21][21] ) );
  OR2X1_RVT U77 ( .A1(\u_div/CryTmp[4][24] ), .A2(\u_div/PartRem[5][24] ), .Y(
        net40598) );
  INVX32_RVT U78 ( .A(\u_div/CryTmp[6][12] ), .Y(n41) );
  IBUFFX4_RVT U79 ( .A(n41), .Y(n42) );
  IBUFFX4_RVT U80 ( .A(\u_div/CryTmp[16][13] ), .Y(n43) );
  IBUFFX4_RVT U81 ( .A(n43), .Y(n44) );
  NBUFFX2_RVT U82 ( .A(net32568), .Y(n45) );
  NBUFFX2_RVT U83 ( .A(net32568), .Y(n46) );
  NBUFFX2_RVT U84 ( .A(net32568), .Y(n47) );
  NBUFFX2_RVT U85 ( .A(net32568), .Y(n48) );
  NBUFFX2_RVT U86 ( .A(net32568), .Y(n49) );
  NBUFFX2_RVT U87 ( .A(net32568), .Y(n50) );
  NBUFFX4_RVT U88 ( .A(net32568), .Y(n51) );
  NBUFFX2_RVT U89 ( .A(net32566), .Y(n52) );
  NBUFFX2_RVT U90 ( .A(net32566), .Y(quotient[15]) );
  NBUFFX2_RVT U91 ( .A(net32566), .Y(n54) );
  NBUFFX2_RVT U92 ( .A(net32566), .Y(n55) );
  NBUFFX2_RVT U93 ( .A(net32566), .Y(n56) );
  NBUFFX2_RVT U94 ( .A(net32566), .Y(n57) );
  NBUFFX4_RVT U95 ( .A(net32566), .Y(n58) );
  IBUFFX4_RVT U96 ( .A(net38340), .Y(n59) );
  IBUFFX16_RVT U97 ( .A(net38340), .Y(net32568) );
  IBUFFX16_RVT U98 ( .A(net38340), .Y(net32566) );
  IBUFFX16_RVT U99 ( .A(net29602), .Y(\u_div/PartRem[9][5] ) );
  MUX21X2_RVT U100 ( .A1(net30184), .A2(net30777), .S0(n194), .Y(n549) );
  INVX4_RVT U101 ( .A(n198), .Y(n194) );
  IBUFFX16_RVT U102 ( .A(n726), .Y(\u_div/PartRem[12][14] ) );
  INVX16_RVT U103 ( .A(n441), .Y(n60) );
  IBUFFX4_RVT U104 ( .A(n60), .Y(n61) );
  IBUFFX8_RVT U105 ( .A(n440), .Y(n441) );
  IBUFFX16_RVT U106 ( .A(\u_div/CryTmp[20][18] ), .Y(n62) );
  IBUFFX2_RVT U107 ( .A(n62), .Y(n63) );
  IBUFFX4_RVT U108 ( .A(\u_div/SumTmp[32][12] ), .Y(n426) );
  INVX4_RVT U109 ( .A(n386), .Y(n64) );
  INVX16_RVT U110 ( .A(n64), .Y(n65) );
  IBUFFX16_RVT U111 ( .A(n378), .Y(n386) );
  IBUFFX4_RVT U112 ( .A(\u_div/CryTmp[4][12] ), .Y(n66) );
  IBUFFX4_RVT U113 ( .A(n66), .Y(n67) );
  IBUFFX16_RVT U114 ( .A(\u_div/SumTmp[2][22] ), .Y(n1143) );
  IBUFFX16_RVT U115 ( .A(n728), .Y(\u_div/PartRem[12][12] ) );
  INVX32_RVT U116 ( .A(\u_div/CryTmp[21][16] ), .Y(n68) );
  IBUFFX16_RVT U117 ( .A(n68), .Y(n69) );
  IBUFFX32_RVT U118 ( .A(\u_div/PartRem[22][12] ), .Y(n70) );
  INVX4_RVT U119 ( .A(n70), .Y(n71) );
  IBUFFX16_RVT U120 ( .A(\u_div/SumTmp[3][19] ), .Y(net30351) );
  IBUFFX16_RVT U121 ( .A(\u_div/CryTmp[23][16] ), .Y(n72) );
  INVX4_RVT U122 ( .A(n72), .Y(n73) );
  INVX8_RVT U123 ( .A(n797), .Y(\u_div/PartRem[6][15] ) );
  MUX21X2_RVT U124 ( .A1(net29666), .A2(net30374), .S0(net45257), .Y(n797) );
  IBUFFX16_RVT U125 ( .A(\u_div/CryTmp[31][12] ), .Y(n438) );
  MUX21X1_RVT U126 ( .A1(net30211), .A2(net29862), .S0(net46343), .Y(net29874)
         );
  INVX8_RVT U127 ( .A(net29862), .Y(\u_div/PartRem[35][10] ) );
  MUX21X2_RVT U128 ( .A1(n1066), .A2(n959), .S0(net50471), .Y(net29862) );
  IBUFFX4_RVT U129 ( .A(\u_div/SumTmp[11][14] ), .Y(net31121) );
  IBUFFX32_RVT U130 ( .A(net31065), .Y(n74) );
  INVX1_RVT U131 ( .A(n74), .Y(n75) );
  IBUFFX16_RVT U132 ( .A(\u_div/SumTmp[4][18] ), .Y(net30352) );
  IBUFFX4_RVT U133 ( .A(\u_div/CryTmp[4][23] ), .Y(n76) );
  INVX2_RVT U134 ( .A(n76), .Y(n77) );
  IBUFFX16_RVT U135 ( .A(net30628), .Y(\u_div/PartRem[17][23] ) );
  INVX2_RVT U136 ( .A(n317), .Y(n318) );
  IBUFFX16_RVT U137 ( .A(\u_div/CryTmp[10][21] ), .Y(n78) );
  INVX4_RVT U138 ( .A(n78), .Y(n79) );
  IBUFFX2_RVT U139 ( .A(\u_div/PartRem[13][10] ), .Y(n80) );
  INVX0_RVT U140 ( .A(n80), .Y(n81) );
  IBUFFX16_RVT U141 ( .A(net30807), .Y(\u_div/PartRem[13][10] ) );
  IBUFFX16_RVT U142 ( .A(\u_div/SumTmp[34][12] ), .Y(n1082) );
  IBUFFX16_RVT U143 ( .A(\u_div/CryTmp[13][10] ), .Y(n82) );
  INVX4_RVT U144 ( .A(n82), .Y(n83) );
  IBUFFX32_RVT U145 ( .A(\u_div/CryTmp[33][14] ), .Y(net31294) );
  IBUFFX16_RVT U146 ( .A(\u_div/SumTmp[25][6] ), .Y(net31011) );
  IBUFFX16_RVT U147 ( .A(net30816), .Y(\u_div/PartRem[13][23] ) );
  MUX21X2_RVT U148 ( .A1(n1193), .A2(n1197), .S0(net42408), .Y(net30816) );
  IBUFFX32_RVT U149 ( .A(\u_div/CryTmp[20][13] ), .Y(n84) );
  IBUFFX4_RVT U150 ( .A(n84), .Y(n85) );
  IBUFFX4_RVT U151 ( .A(net29898), .Y(\u_div/PartRem[32][1] ) );
  NBUFFX8_RVT U152 ( .A(net32550), .Y(quotient[12]) );
  NBUFFX32_RVT U153 ( .A(net32550), .Y(n87) );
  INVX0_RVT U154 ( .A(net38337), .Y(net32550) );
  INVX1_RVT U155 ( .A(\u_div/CryTmp[21][9] ), .Y(n181) );
  IBUFFX16_RVT U156 ( .A(\u_div/CryTmp[5][15] ), .Y(n88) );
  INVX4_RVT U157 ( .A(n88), .Y(n89) );
  INVX1_RVT U158 ( .A(\u_div/PartRem[28][13] ), .Y(net49678) );
  INVX4_RVT U159 ( .A(net31056), .Y(n90) );
  IBUFFX16_RVT U160 ( .A(n90), .Y(n91) );
  IBUFFX16_RVT U161 ( .A(\u_div/CryTmp[23][8] ), .Y(n92) );
  INVX4_RVT U162 ( .A(n92), .Y(n93) );
  IBUFFX16_RVT U163 ( .A(\u_div/CryTmp[45][2] ), .Y(n94) );
  INVX4_RVT U164 ( .A(n94), .Y(n95) );
  IBUFFX4_RVT U165 ( .A(\u_div/CryTmp[16][23] ), .Y(n96) );
  INVX4_RVT U166 ( .A(n96), .Y(n97) );
  IBUFFX4_RVT U167 ( .A(\u_div/PartRem[12][13] ), .Y(n98) );
  IBUFFX16_RVT U168 ( .A(n98), .Y(n99) );
  IBUFFX16_RVT U169 ( .A(n727), .Y(\u_div/PartRem[12][13] ) );
  IBUFFX16_RVT U170 ( .A(\u_div/CryTmp[15][16] ), .Y(n100) );
  INVX4_RVT U171 ( .A(n100), .Y(n101) );
  IBUFFX32_RVT U172 ( .A(n767), .Y(n102) );
  INVX1_RVT U173 ( .A(n102), .Y(n103) );
  IBUFFX16_RVT U174 ( .A(net30863), .Y(\u_div/PartRem[12][23] ) );
  IBUFFX4_RVT U175 ( .A(\u_div/CryTmp[11][23] ), .Y(n104) );
  INVX2_RVT U176 ( .A(n104), .Y(n105) );
  IBUFFX4_RVT U177 ( .A(n444), .Y(n445) );
  INVX32_RVT U178 ( .A(\u_div/CryTmp[28][13] ), .Y(n106) );
  IBUFFX16_RVT U179 ( .A(n106), .Y(n107) );
  IBUFFX16_RVT U180 ( .A(\u_div/CryTmp[11][10] ), .Y(n108) );
  INVX4_RVT U181 ( .A(n108), .Y(n109) );
  IBUFFX16_RVT U182 ( .A(\u_div/CryTmp[20][17] ), .Y(n110) );
  INVX4_RVT U183 ( .A(n110), .Y(n111) );
  INVX2_RVT U184 ( .A(n901), .Y(n902) );
  INVX4_RVT U185 ( .A(net48385), .Y(net47978) );
  IBUFFX16_RVT U186 ( .A(\u_div/SumTmp[14][22] ), .Y(n1195) );
  MUX21X2_RVT U187 ( .A1(net30528), .A2(net31144), .S0(net32580), .Y(n646) );
  IBUFFX16_RVT U188 ( .A(net30528), .Y(\u_div/PartRem[18][7] ) );
  MUX21X2_RVT U189 ( .A1(n600), .A2(net31145), .S0(net45678), .Y(net30528) );
  INVX8_RVT U190 ( .A(n115), .Y(net48384) );
  INVX32_RVT U191 ( .A(\u_div/CryTmp[9][18] ), .Y(n112) );
  IBUFFX16_RVT U192 ( .A(n112), .Y(n113) );
  IBUFFX4_RVT U193 ( .A(net32596), .Y(n114) );
  INVX32_RVT U194 ( .A(n114), .Y(n115) );
  IBUFFX16_RVT U195 ( .A(\u_div/SumTmp[43][3] ), .Y(n357) );
  IBUFFX16_RVT U196 ( .A(\u_div/CryTmp[14][18] ), .Y(n116) );
  INVX4_RVT U197 ( .A(n116), .Y(n117) );
  AND3X4_RVT U198 ( .A1(net47690), .A2(net31938), .A3(\u_div/CryTmp[29][18] ), 
        .Y(net47679) );
  IBUFFX4_RVT U199 ( .A(\u_div/CryTmp[8][5] ), .Y(n118) );
  IBUFFX4_RVT U200 ( .A(n118), .Y(n119) );
  IBUFFX4_RVT U201 ( .A(n1230), .Y(n120) );
  INVX2_RVT U202 ( .A(n120), .Y(n121) );
  IBUFFX8_RVT U203 ( .A(\u_div/PartRem[21][12] ), .Y(n122) );
  IBUFFX4_RVT U204 ( .A(n122), .Y(n123) );
  IBUFFX4_RVT U205 ( .A(net30277), .Y(\u_div/PartRem[20][16] ) );
  IBUFFX4_RVT U206 ( .A(\u_div/PartRem[5][19] ), .Y(n124) );
  INVX2_RVT U207 ( .A(n124), .Y(n125) );
  INVX0_RVT U208 ( .A(n812), .Y(\u_div/PartRem[5][19] ) );
  IBUFFX4_RVT U209 ( .A(\u_div/CryTmp[13][23] ), .Y(n126) );
  IBUFFX4_RVT U210 ( .A(n126), .Y(n127) );
  IBUFFX16_RVT U211 ( .A(\u_div/SumTmp[3][13] ), .Y(net30411) );
  INVX0_RVT U212 ( .A(n854), .Y(n128) );
  INVX1_RVT U213 ( .A(n854), .Y(quotient[5]) );
  OR2X2_RVT U214 ( .A1(\u_div/PartRem[6][24] ), .A2(\u_div/CryTmp[5][24] ), 
        .Y(net49616) );
  INVX2_RVT U215 ( .A(net45654), .Y(net49611) );
  INVX2_RVT U216 ( .A(net49612), .Y(net49625) );
  INVX2_RVT U217 ( .A(net49626), .Y(net32506) );
  INVX2_RVT U218 ( .A(n854), .Y(net44755) );
  IBUFFX16_RVT U219 ( .A(net49616), .Y(net45654) );
  IBUFFX4_RVT U220 ( .A(net49611), .Y(net49612) );
  IBUFFX4_RVT U221 ( .A(net49625), .Y(net49626) );
  IBUFFX4_RVT U222 ( .A(net32506), .Y(n854) );
  IBUFFX4_RVT U223 ( .A(\u_div/CryTmp[16][18] ), .Y(n130) );
  IBUFFX4_RVT U224 ( .A(n130), .Y(n131) );
  IBUFFX16_RVT U225 ( .A(\u_div/SumTmp[28][15] ), .Y(n1126) );
  IBUFFX16_RVT U226 ( .A(\u_div/CryTmp[18][23] ), .Y(n132) );
  INVX4_RVT U227 ( .A(n132), .Y(n133) );
  IBUFFX16_RVT U228 ( .A(\u_div/CryTmp[23][22] ), .Y(n134) );
  INVX4_RVT U229 ( .A(n134), .Y(n135) );
  IBUFFX16_RVT U230 ( .A(\u_div/CryTmp[18][8] ), .Y(n136) );
  INVX4_RVT U231 ( .A(n136), .Y(n137) );
  IBUFFX16_RVT U232 ( .A(net30006), .Y(\u_div/PartRem[26][7] ) );
  IBUFFX16_RVT U233 ( .A(\u_div/SumTmp[25][21] ), .Y(net30079) );
  INVX32_RVT U234 ( .A(\u_div/CryTmp[9][16] ), .Y(n138) );
  IBUFFX16_RVT U235 ( .A(n138), .Y(n139) );
  NOR3X0_RVT U236 ( .A1(net31872), .A2(net31315), .A3(n484), .Y(n140) );
  NOR3X0_RVT U237 ( .A1(net31872), .A2(net31315), .A3(n484), .Y(n141) );
  IBUFFX4_RVT U238 ( .A(n140), .Y(n142) );
  IBUFFX4_RVT U239 ( .A(n142), .Y(n143) );
  IBUFFX4_RVT U240 ( .A(n142), .Y(n144) );
  IBUFFX4_RVT U241 ( .A(n142), .Y(n145) );
  IBUFFX16_RVT U242 ( .A(n141), .Y(n146) );
  IBUFFX4_RVT U243 ( .A(n146), .Y(quotient[26]) );
  IBUFFX4_RVT U244 ( .A(n146), .Y(n148) );
  INVX4_RVT U245 ( .A(n146), .Y(n149) );
  IBUFFX16_RVT U246 ( .A(net37567), .Y(n150) );
  IBUFFX4_RVT U247 ( .A(n150), .Y(n151) );
  IBUFFX4_RVT U248 ( .A(n150), .Y(n152) );
  INVX4_RVT U249 ( .A(n150), .Y(n153) );
  NOR3X0_RVT U250 ( .A1(net31872), .A2(net31315), .A3(n484), .Y(net37567) );
  IBUFFX16_RVT U251 ( .A(\u_div/SumTmp[3][12] ), .Y(net30421) );
  IBUFFX16_RVT U252 ( .A(\u_div/CryTmp[16][7] ), .Y(n154) );
  INVX4_RVT U253 ( .A(n154), .Y(n155) );
  MUX21X2_RVT U254 ( .A1(net30279), .A2(net30955), .S0(net32590), .Y(n611) );
  IBUFFX16_RVT U255 ( .A(net30279), .Y(\u_div/PartRem[20][14] ) );
  IBUFFX4_RVT U256 ( .A(net32578), .Y(n156) );
  IBUFFX4_RVT U257 ( .A(n156), .Y(n157) );
  INVX4_RVT U258 ( .A(n156), .Y(n158) );
  IBUFFX32_RVT U259 ( .A(\u_div/CryTmp[20][12] ), .Y(n159) );
  IBUFFX4_RVT U260 ( .A(n159), .Y(n160) );
  INVX4_RVT U261 ( .A(n629), .Y(n161) );
  IBUFFX8_RVT U262 ( .A(n161), .Y(n162) );
  IBUFFX4_RVT U263 ( .A(n165), .Y(n163) );
  INVX1_RVT U264 ( .A(n163), .Y(n164) );
  IBUFFX16_RVT U265 ( .A(\u_div/CryTmp[24][21] ), .Y(n165) );
  IBUFFX4_RVT U266 ( .A(n164), .Y(n166) );
  INVX32_RVT U267 ( .A(\u_div/PartRem[42][2] ), .Y(n167) );
  IBUFFX4_RVT U268 ( .A(n167), .Y(n168) );
  INVX2_RVT U269 ( .A(n576), .Y(n169) );
  IBUFFX4_RVT U270 ( .A(n169), .Y(n170) );
  NBUFFX8_RVT U271 ( .A(net47716), .Y(n171) );
  NBUFFX8_RVT U272 ( .A(net47716), .Y(n172) );
  NBUFFX8_RVT U273 ( .A(net47716), .Y(quotient[39]) );
  IBUFFX16_RVT U274 ( .A(\u_div/CryTmp[20][15] ), .Y(n174) );
  INVX4_RVT U275 ( .A(n174), .Y(n175) );
  OR2X1_RVT U276 ( .A1(\u_div/CryTmp[4][24] ), .A2(\u_div/PartRem[5][24] ), 
        .Y(n176) );
  IBUFFX4_RVT U277 ( .A(net50726), .Y(net50727) );
  NAND2X4_RVT U278 ( .A1(n33), .A2(\u_div/CryTmp[22][16] ), .Y(n583) );
  IBUFFX16_RVT U279 ( .A(net30124), .Y(\u_div/PartRem[23][16] ) );
  IBUFFX4_RVT U280 ( .A(\u_div/CryTmp[26][13] ), .Y(n177) );
  INVX2_RVT U281 ( .A(n177), .Y(n178) );
  IBUFFX4_RVT U282 ( .A(\u_div/PartRem[25][9] ), .Y(n179) );
  INVX2_RVT U283 ( .A(n179), .Y(n180) );
  IBUFFX4_RVT U284 ( .A(n181), .Y(n182) );
  IBUFFX16_RVT U285 ( .A(\u_div/CryTmp[35][11] ), .Y(n960) );
  NBUFFX16_RVT U286 ( .A(net32616), .Y(quotient[23]) );
  INVX4_RVT U287 ( .A(n558), .Y(net32616) );
  IBUFFX16_RVT U288 ( .A(\u_div/SumTmp[12][18] ), .Y(net31021) );
  NOR2X2_RVT U289 ( .A1(\u_div/CryTmp[19][24] ), .A2(\u_div/PartRem[20][24] ), 
        .Y(net38344) );
  IBUFFX16_RVT U290 ( .A(\u_div/CryTmp[2][19] ), .Y(n901) );
  IBUFFX16_RVT U291 ( .A(\u_div/CryTmp[9][14] ), .Y(n184) );
  INVX4_RVT U292 ( .A(n184), .Y(n185) );
  IBUFFX32_RVT U293 ( .A(n185), .Y(n186) );
  IBUFFX4_RVT U294 ( .A(n186), .Y(n187) );
  INVX2_RVT U295 ( .A(net37585), .Y(net50470) );
  IBUFFX4_RVT U296 ( .A(n742), .Y(n743) );
  IBUFFX4_RVT U297 ( .A(net30762), .Y(\u_div/PartRem[13][8] ) );
  INVX2_RVT U298 ( .A(n643), .Y(n644) );
  IBUFFX4_RVT U299 ( .A(\u_div/SumTmp[3][11] ), .Y(net30431) );
  INVX2_RVT U300 ( .A(n1051), .Y(\u_div/PartRem[3][12] ) );
  MUX21X2_RVT U301 ( .A1(net30806), .A2(net31155), .S0(quotient[12]), .Y(n728)
         );
  IBUFFX16_RVT U302 ( .A(net30806), .Y(\u_div/PartRem[13][11] ) );
  MUX21X2_RVT U303 ( .A1(n714), .A2(net31156), .S0(net32554), .Y(net30806) );
  MUX21X2_RVT U304 ( .A1(\u_div/PartRem[22][23] ), .A2(\u_div/SumTmp[21][23] ), 
        .S0(quotient[21]), .Y(\u_div/PartRem[21][24] ) );
  IBUFFX2_RVT U305 ( .A(n197), .Y(quotient[21]) );
  IBUFFX4_RVT U306 ( .A(\u_div/PartRem[14][7] ), .Y(n188) );
  INVX4_RVT U307 ( .A(n188), .Y(n189) );
  NOR2X4_RVT U308 ( .A1(net31814), .A2(net31320), .Y(net47709) );
  IBUFFX32_RVT U309 ( .A(\u_div/CryTmp[24][23] ), .Y(net31320) );
  IBUFFX4_RVT U310 ( .A(\u_div/CryTmp[11][24] ), .Y(net46895) );
  IBUFFX16_RVT U311 ( .A(net38342), .Y(n190) );
  IBUFFX4_RVT U312 ( .A(net38342), .Y(n191) );
  IBUFFX4_RVT U313 ( .A(n196), .Y(n192) );
  IBUFFX4_RVT U314 ( .A(n197), .Y(n193) );
  IBUFFX32_RVT U315 ( .A(n198), .Y(n195) );
  INVX1_RVT U316 ( .A(n190), .Y(n196) );
  INVX1_RVT U317 ( .A(n190), .Y(n197) );
  INVX1_RVT U318 ( .A(n190), .Y(n198) );
  INVX1_RVT U319 ( .A(n196), .Y(n199) );
  INVX1_RVT U320 ( .A(n196), .Y(n200) );
  INVX1_RVT U321 ( .A(n196), .Y(n201) );
  INVX1_RVT U322 ( .A(n196), .Y(n202) );
  INVX1_RVT U323 ( .A(n197), .Y(n203) );
  INVX1_RVT U324 ( .A(n197), .Y(n204) );
  INVX1_RVT U325 ( .A(n197), .Y(n205) );
  INVX1_RVT U326 ( .A(n198), .Y(n207) );
  INVX1_RVT U327 ( .A(n198), .Y(n208) );
  INVX1_RVT U328 ( .A(n198), .Y(n209) );
  INVX1_RVT U329 ( .A(n198), .Y(n210) );
  IBUFFX16_RVT U330 ( .A(\u_div/SumTmp[37][4] ), .Y(n1182) );
  IBUFFX16_RVT U331 ( .A(\u_div/CryTmp[3][6] ), .Y(n843) );
  INVX4_RVT U332 ( .A(n917), .Y(n918) );
  IBUFFX16_RVT U333 ( .A(\u_div/CryTmp[2][12] ), .Y(n917) );
  INVX1_RVT U334 ( .A(net38344), .Y(n211) );
  INVX8_RVT U335 ( .A(net38344), .Y(n212) );
  INVX4_RVT U336 ( .A(net42365), .Y(net32590) );
  IBUFFX4_RVT U337 ( .A(n866), .Y(n868) );
  IBUFFX16_RVT U338 ( .A(\u_div/CryTmp[22][15] ), .Y(n213) );
  INVX4_RVT U339 ( .A(n213), .Y(n214) );
  IBUFFX16_RVT U340 ( .A(\u_div/CryTmp[5][22] ), .Y(n215) );
  INVX4_RVT U341 ( .A(n215), .Y(n216) );
  IBUFFX16_RVT U342 ( .A(\u_div/CryTmp[41][4] ), .Y(n217) );
  INVX4_RVT U343 ( .A(n217), .Y(n218) );
  OR2X2_RVT U344 ( .A1(\u_div/PartRem[1][24] ), .A2(\u_div/CryTmp[0][24] ), 
        .Y(quotient[0]) );
  IBUFFX16_RVT U345 ( .A(\u_div/CryTmp[0][23] ), .Y(n219) );
  IBUFFX16_RVT U346 ( .A(n219), .Y(n220) );
  IBUFFX4_RVT U347 ( .A(\u_div/CryTmp[1][16] ), .Y(n221) );
  IBUFFX4_RVT U348 ( .A(n221), .Y(n222) );
  IBUFFX16_RVT U349 ( .A(net29603), .Y(\u_div/PartRem[9][4] ) );
  INVX4_RVT U350 ( .A(n511), .Y(n223) );
  IBUFFX16_RVT U351 ( .A(n223), .Y(n224) );
  IBUFFX4_RVT U352 ( .A(\u_div/CryTmp[1][22] ), .Y(n225) );
  IBUFFX4_RVT U353 ( .A(n225), .Y(n226) );
  IBUFFX4_RVT U354 ( .A(\u_div/CryTmp[21][21] ), .Y(n227) );
  IBUFFX4_RVT U355 ( .A(n227), .Y(n228) );
  INVX32_RVT U356 ( .A(\u_div/CryTmp[32][13] ), .Y(n229) );
  IBUFFX16_RVT U357 ( .A(n229), .Y(n230) );
  INVX2_RVT U358 ( .A(n625), .Y(n626) );
  INVX2_RVT U359 ( .A(net31243), .Y(n231) );
  IBUFFX4_RVT U360 ( .A(n231), .Y(n232) );
  IBUFFX4_RVT U361 ( .A(\u_div/PartRem[35][1] ), .Y(n233) );
  INVX4_RVT U362 ( .A(n233), .Y(n234) );
  INVX1_RVT U363 ( .A(n398), .Y(\u_div/PartRem[35][1] ) );
  IBUFFX4_RVT U364 ( .A(n438), .Y(n439) );
  INVX2_RVT U365 ( .A(n679), .Y(n680) );
  IBUFFX16_RVT U366 ( .A(\u_div/CryTmp[27][9] ), .Y(n235) );
  INVX4_RVT U367 ( .A(n235), .Y(n236) );
  INVX4_RVT U368 ( .A(n631), .Y(n237) );
  IBUFFX8_RVT U369 ( .A(n237), .Y(n238) );
  INVX4_RVT U370 ( .A(net31303), .Y(n239) );
  IBUFFX16_RVT U371 ( .A(n239), .Y(n240) );
  INVX4_RVT U372 ( .A(n563), .Y(n241) );
  IBUFFX8_RVT U373 ( .A(n241), .Y(n242) );
  IBUFFX16_RVT U374 ( .A(n847), .Y(n867) );
  INVX32_RVT U375 ( .A(\u_div/CryTmp[3][23] ), .Y(n847) );
  INVX4_RVT U376 ( .A(n862), .Y(n863) );
  IBUFFX16_RVT U377 ( .A(\u_div/CryTmp[3][12] ), .Y(n862) );
  IBUFFX4_RVT U378 ( .A(\u_div/PartRem[9][3] ), .Y(n243) );
  IBUFFX4_RVT U379 ( .A(n243), .Y(n244) );
  IBUFFX16_RVT U380 ( .A(net29604), .Y(\u_div/PartRem[9][3] ) );
  IBUFFX32_RVT U381 ( .A(n310), .Y(n245) );
  IBUFFX4_RVT U382 ( .A(n245), .Y(n246) );
  IBUFFX16_RVT U383 ( .A(\u_div/CryTmp[29][10] ), .Y(n247) );
  INVX4_RVT U384 ( .A(n247), .Y(n248) );
  IBUFFX16_RVT U385 ( .A(\u_div/CryTmp[26][10] ), .Y(n249) );
  INVX4_RVT U386 ( .A(n249), .Y(n250) );
  IBUFFX16_RVT U387 ( .A(\u_div/CryTmp[4][6] ), .Y(n251) );
  INVX4_RVT U388 ( .A(n251), .Y(n252) );
  IBUFFX16_RVT U389 ( .A(\u_div/CryTmp[32][8] ), .Y(n253) );
  INVX2_RVT U390 ( .A(n253), .Y(n254) );
  MUX21X2_RVT U391 ( .A1(n780), .A2(net30290), .S0(net46768), .Y(n784) );
  INVX32_RVT U392 ( .A(n780), .Y(\u_div/PartRem[8][2] ) );
  MUX21X2_RVT U393 ( .A1(net29609), .A2(net30291), .S0(net40719), .Y(n780) );
  IBUFFX16_RVT U394 ( .A(\u_div/CryTmp[17][2] ), .Y(n255) );
  INVX4_RVT U395 ( .A(n255), .Y(n256) );
  IBUFFX16_RVT U396 ( .A(\u_div/CryTmp[3][4] ), .Y(n257) );
  INVX4_RVT U397 ( .A(n257), .Y(n258) );
  IBUFFX32_RVT U398 ( .A(net29636), .Y(n259) );
  IBUFFX4_RVT U399 ( .A(n259), .Y(n260) );
  MUX21X2_RVT U400 ( .A1(net29612), .A2(net29944), .S0(net40719), .Y(net29636)
         );
  IBUFFX4_RVT U401 ( .A(\u_div/CryTmp[7][17] ), .Y(n261) );
  IBUFFX4_RVT U402 ( .A(n261), .Y(n262) );
  IBUFFX4_RVT U403 ( .A(\u_div/CryTmp[7][8] ), .Y(n263) );
  IBUFFX4_RVT U404 ( .A(n263), .Y(n264) );
  IBUFFX4_RVT U405 ( .A(\u_div/CryTmp[7][12] ), .Y(n265) );
  IBUFFX4_RVT U406 ( .A(n265), .Y(n266) );
  IBUFFX16_RVT U407 ( .A(\u_div/CryTmp[4][19] ), .Y(n267) );
  INVX4_RVT U408 ( .A(n267), .Y(n268) );
  IBUFFX16_RVT U409 ( .A(\u_div/CryTmp[21][15] ), .Y(n269) );
  INVX4_RVT U410 ( .A(n269), .Y(n270) );
  IBUFFX4_RVT U411 ( .A(\u_div/CryTmp[0][17] ), .Y(n271) );
  IBUFFX4_RVT U412 ( .A(n271), .Y(n272) );
  IBUFFX32_RVT U413 ( .A(n887), .Y(n273) );
  INVX8_RVT U414 ( .A(n273), .Y(n274) );
  IBUFFX16_RVT U415 ( .A(\u_div/CryTmp[3][2] ), .Y(n275) );
  INVX4_RVT U416 ( .A(n275), .Y(n276) );
  IBUFFX4_RVT U417 ( .A(n392), .Y(n277) );
  IBUFFX4_RVT U418 ( .A(n277), .Y(n278) );
  MUX21X1_RVT U419 ( .A1(net29841), .A2(net30260), .S0(net50471), .Y(n392) );
  IBUFFX4_RVT U420 ( .A(net30843), .Y(n279) );
  IBUFFX4_RVT U421 ( .A(n279), .Y(n280) );
  MUX21X1_RVT U422 ( .A1(net30798), .A2(net30998), .S0(net32548), .Y(net30843)
         );
  INVX32_RVT U423 ( .A(n280), .Y(\u_div/PartRem[12][20] ) );
  NOR2X4_RVT U424 ( .A1(\u_div/PartRem[9][24] ), .A2(\u_div/CryTmp[8][24] ), 
        .Y(net47729) );
  INVX4_RVT U425 ( .A(net40717), .Y(net40719) );
  IBUFFX4_RVT U426 ( .A(net40717), .Y(net40721) );
  IBUFFX4_RVT U427 ( .A(net40717), .Y(net40720) );
  IBUFFX4_RVT U428 ( .A(net40717), .Y(net40718) );
  MUX21X1_RVT U429 ( .A1(n419), .A2(n426), .S0(n435), .Y(net29901) );
  INVX1_RVT U430 ( .A(n335), .Y(\u_div/PartRem[43][1] ) );
  IBUFFX4_RVT U431 ( .A(\u_div/SumTmp[33][12] ), .Y(net30150) );
  MUX21X1_RVT U432 ( .A1(net30053), .A2(net31115), .S0(quotient[23]), .Y(
        net30074) );
  MUX21X1_RVT U433 ( .A1(net30021), .A2(net30685), .S0(quotient[25]), .Y(n499)
         );
  INVX1_RVT U434 ( .A(\u_div/SumTmp[33][8] ), .Y(net30549) );
  MUX21X1_RVT U435 ( .A1(n692), .A2(n733), .S0(net32560), .Y(n709) );
  IBUFFX4_RVT U436 ( .A(net29852), .Y(\u_div/PartRem[35][8] ) );
  INVX1_RVT U437 ( .A(\u_div/CryTmp[21][20] ), .Y(n1004) );
  INVX1_RVT U438 ( .A(n958), .Y(n959) );
  INVX0_RVT U439 ( .A(n1122), .Y(n958) );
  MUX21X1_RVT U440 ( .A1(n334), .A2(net30219), .S0(net37556), .Y(n387) );
  INVX1_RVT U441 ( .A(\u_div/SumTmp[31][14] ), .Y(net30148) );
  MUX21X1_RVT U442 ( .A1(net29885), .A2(net30086), .S0(net50050), .Y(net29899)
         );
  MUX21X1_RVT U443 ( .A1(n533), .A2(n557), .S0(net32608), .Y(net30134) );
  MUX21X1_RVT U444 ( .A1(net31642), .A2(net37254), .S0(net50049), .Y(net29898)
         );
  INVX0_RVT U445 ( .A(n702), .Y(\u_div/PartRem[14][5] ) );
  INVX1_RVT U446 ( .A(net29913), .Y(\u_div/PartRem[31][1] ) );
  MUX21X1_RVT U447 ( .A1(n417), .A2(net30968), .S0(net50050), .Y(net29897) );
  MUX21X1_RVT U448 ( .A1(n416), .A2(net30884), .S0(net50049), .Y(net29896) );
  MUX21X1_RVT U449 ( .A1(n541), .A2(net31073), .S0(net44969), .Y(net30237) );
  MUX21X1_RVT U450 ( .A1(net29968), .A2(net30963), .S0(net41415), .Y(net29986)
         );
  MUX21X1_RVT U451 ( .A1(net30004), .A2(net30877), .S0(quotient[25]), .Y(
        net41435) );
  INVX1_RVT U452 ( .A(net29966), .Y(\u_div/PartRem[28][8] ) );
  INVX1_RVT U453 ( .A(\u_div/PartRem[20][14] ), .Y(n587) );
  MUX21X1_RVT U454 ( .A1(net45295), .A2(net30732), .S0(net47709), .Y(net30064)
         );
  MUX21X1_RVT U455 ( .A1(net30357), .A2(net30358), .S0(net32530), .Y(net29615)
         );
  INVX1_RVT U456 ( .A(n515), .Y(n516) );
  INVX1_RVT U457 ( .A(\u_div/CryTmp[24][14] ), .Y(n515) );
  MUX21X1_RVT U458 ( .A1(net30277), .A2(net30823), .S0(n212), .Y(n609) );
  MUX21X1_RVT U459 ( .A1(net30123), .A2(net30634), .S0(net32610), .Y(net30181)
         );
  INVX1_RVT U460 ( .A(\u_div/SumTmp[36][5] ), .Y(n1181) );
  MUX21X1_RVT U461 ( .A1(net29817), .A2(net30506), .S0(net37581), .Y(n1056) );
  INVX1_RVT U462 ( .A(net30845), .Y(\u_div/PartRem[12][19] ) );
  MUX21X1_RVT U463 ( .A1(n708), .A2(net30975), .S0(net42408), .Y(net30796) );
  INVX1_RVT U464 ( .A(net30017), .Y(\u_div/PartRem[26][17] ) );
  MUX21X1_RVT U465 ( .A1(n335), .A2(net30267), .S0(net37556), .Y(n338) );
  INVX1_RVT U466 ( .A(net29977), .Y(\u_div/PartRem[28][16] ) );
  INVX0_RVT U467 ( .A(net37563), .Y(net46343) );
  IBUFFX4_RVT U468 ( .A(\u_div/SumTmp[34][10] ), .Y(net30211) );
  INVX1_RVT U469 ( .A(n334), .Y(\u_div/PartRem[43][2] ) );
  IBUFFX4_RVT U470 ( .A(\u_div/SumTmp[35][10] ), .Y(n1105) );
  INVX1_RVT U471 ( .A(\u_div/SumTmp[41][5] ), .Y(n355) );
  INVX1_RVT U472 ( .A(n1119), .Y(\u_div/PartRem[22][22] ) );
  MUX21X1_RVT U473 ( .A1(\u_div/PartRem[25][22] ), .A2(\u_div/SumTmp[24][22] ), 
        .S0(net47709), .Y(n559) );
  INVX1_RVT U474 ( .A(\u_div/SumTmp[36][10] ), .Y(n1084) );
  MUX21X1_RVT U475 ( .A1(n607), .A2(net31212), .S0(n635), .Y(net30533) );
  INVX1_RVT U476 ( .A(n570), .Y(n571) );
  INVX1_RVT U477 ( .A(\u_div/CryTmp[20][6] ), .Y(n570) );
  MUX21X1_RVT U478 ( .A1(net30891), .A2(net30944), .S0(net32536), .Y(net30467)
         );
  NBUFFX4_RVT U479 ( .A(net31016), .Y(net52534) );
  INVX1_RVT U480 ( .A(\u_div/SumTmp[30][1] ), .Y(net31016) );
  INVX1_RVT U481 ( .A(n701), .Y(\u_div/PartRem[14][6] ) );
  INVX0_RVT U482 ( .A(n103), .Y(n768) );
  INVX0_RVT U483 ( .A(n224), .Y(n512) );
  MUX21X1_RVT U484 ( .A1(net30004), .A2(net30877), .S0(quotient[25]), .Y(n501)
         );
  INVX2_RVT U485 ( .A(n453), .Y(n454) );
  MUX21X1_RVT U486 ( .A1(net29895), .A2(net30835), .S0(net40084), .Y(net29909)
         );
  MUX21X1_RVT U487 ( .A1(net30068), .A2(net30959), .S0(quotient[23]), .Y(n1102) );
  IBUFFX4_RVT U488 ( .A(\u_div/SumTmp[13][10] ), .Y(net31156) );
  INVX1_RVT U489 ( .A(\u_div/SumTmp[27][9] ), .Y(net30783) );
  INVX1_RVT U490 ( .A(\u_div/CryTmp[8][11] ), .Y(n773) );
  MUX21X1_RVT U491 ( .A1(net29907), .A2(net30738), .S0(net37577), .Y(n457) );
  INVX1_RVT U492 ( .A(\u_div/SumTmp[20][14] ), .Y(net30872) );
  INVX0_RVT U493 ( .A(n305), .Y(n306) );
  INVX1_RVT U494 ( .A(net30896), .Y(\u_div/PartRem[11][15] ) );
  IBUFFX4_RVT U495 ( .A(\u_div/CryTmp[10][15] ), .Y(n305) );
  MUX21X1_RVT U496 ( .A1(n499), .A2(net30684), .S0(net47709), .Y(net30063) );
  INVX1_RVT U497 ( .A(n496), .Y(n494) );
  INVX1_RVT U498 ( .A(n495), .Y(n496) );
  NAND2X1_RVT U499 ( .A1(\u_div/PartRem[23][15] ), .A2(n214), .Y(net49310) );
  INVX1_RVT U500 ( .A(n589), .Y(n590) );
  MUX21X1_RVT U501 ( .A1(net30040), .A2(net30588), .S0(net47709), .Y(n531) );
  INVX1_RVT U502 ( .A(net29819), .Y(\u_div/PartRem[39][2] ) );
  INVX0_RVT U503 ( .A(n943), .Y(n944) );
  INVX1_RVT U504 ( .A(n1021), .Y(\u_div/PartRem[8][16] ) );
  INVX0_RVT U505 ( .A(n678), .Y(\u_div/PartRem[16][17] ) );
  INVX1_RVT U506 ( .A(n401), .Y(\u_div/PartRem[34][7] ) );
  MUX21X1_RVT U507 ( .A1(n345), .A2(net30556), .S0(net50177), .Y(n349) );
  INVX1_RVT U508 ( .A(net50176), .Y(net50177) );
  INVX1_RVT U509 ( .A(net49212), .Y(net50176) );
  INVX1_RVT U510 ( .A(\u_div/SumTmp[31][12] ), .Y(net30256) );
  MUX21X1_RVT U511 ( .A1(net31466), .A2(net37224), .S0(quotient[43]), .Y(n335)
         );
  MUX21X1_RVT U512 ( .A1(n761), .A2(net29738), .S0(net40720), .Y(net29633) );
  INVX1_RVT U513 ( .A(n937), .Y(n938) );
  MUX21X1_RVT U514 ( .A1(n593), .A2(net30632), .S0(net32598), .Y(n595) );
  MUX21X1_RVT U515 ( .A1(n278), .A2(n446), .S0(net37563), .Y(n408) );
  INVX1_RVT U516 ( .A(\u_div/SumTmp[34][9] ), .Y(n446) );
  MUX21X1_RVT U517 ( .A1(net30845), .A2(net31020), .S0(net32542), .Y(net30890)
         );
  MUX21X1_RVT U518 ( .A1(n280), .A2(net30997), .S0(net32542), .Y(net30889) );
  MUX21X1_RVT U519 ( .A1(n373), .A2(n374), .S0(quotient[44]), .Y(n331) );
  INVX1_RVT U520 ( .A(n775), .Y(\u_div/PartRem[9][21] ) );
  MUX21X1_RVT U521 ( .A1(n706), .A2(n730), .S0(net42408), .Y(net30795) );
  INVX1_RVT U522 ( .A(net52401), .Y(net52402) );
  INVX1_RVT U523 ( .A(net30654), .Y(\u_div/PartRem[16][21] ) );
  INVX2_RVT U524 ( .A(n26), .Y(n292) );
  INVX1_RVT U525 ( .A(net30015), .Y(\u_div/PartRem[26][19] ) );
  INVX1_RVT U526 ( .A(net29916), .Y(\u_div/PartRem[31][14] ) );
  INVX1_RVT U527 ( .A(n418), .Y(\u_div/PartRem[33][13] ) );
  INVX1_RVT U528 ( .A(net49211), .Y(n385) );
  INVX4_RVT U529 ( .A(n170), .Y(n577) );
  INVX1_RVT U530 ( .A(net38346), .Y(net32578) );
  IBUFFX4_RVT U531 ( .A(net29975), .Y(\u_div/PartRem[28][18] ) );
  INVX1_RVT U532 ( .A(n332), .Y(\u_div/PartRem[43][4] ) );
  INVX1_RVT U533 ( .A(b[13]), .Y(net32078) );
  INVX1_RVT U534 ( .A(b[3]), .Y(net32354) );
  INVX1_RVT U535 ( .A(net31974), .Y(net31972) );
  INVX0_RVT U536 ( .A(\u_div/PartRem[28][19] ), .Y(net44394) );
  INVX1_RVT U537 ( .A(net29974), .Y(\u_div/PartRem[28][19] ) );
  INVX1_RVT U538 ( .A(net32242), .Y(net32234) );
  INVX1_RVT U539 ( .A(n960), .Y(n961) );
  INVX1_RVT U540 ( .A(net41045), .Y(net30036) );
  INVX1_RVT U541 ( .A(n604), .Y(\u_div/PartRem[19][2] ) );
  INVX1_RVT U542 ( .A(\u_div/SumTmp[24][3] ), .Y(net31097) );
  MUX21X1_RVT U543 ( .A1(net30627), .A2(net30916), .S0(n47), .Y(n687) );
  INVX2_RVT U544 ( .A(n289), .Y(n290) );
  INVX1_RVT U545 ( .A(n651), .Y(\u_div/PartRem[17][3] ) );
  INVX1_RVT U546 ( .A(\u_div/CryTmp[16][3] ), .Y(n289) );
  INVX0_RVT U547 ( .A(net46688), .Y(net30135) );
  INVX1_RVT U548 ( .A(n503), .Y(n505) );
  INVX1_RVT U549 ( .A(\u_div/CryTmp[25][4] ), .Y(n503) );
  INVX1_RVT U550 ( .A(\u_div/SumTmp[26][3] ), .Y(net31057) );
  INVX1_RVT U551 ( .A(net30626), .Y(\u_div/PartRem[16][3] ) );
  INVX1_RVT U552 ( .A(\u_div/SumTmp[21][6] ), .Y(net31094) );
  MUX21X1_RVT U553 ( .A1(net31674), .A2(net37261), .S0(net37577), .Y(n464) );
  INVX2_RVT U554 ( .A(n487), .Y(n488) );
  INVX1_RVT U555 ( .A(net29971), .Y(\u_div/PartRem[28][3] ) );
  INVX1_RVT U556 ( .A(\u_div/SumTmp[26][5] ), .Y(net31012) );
  INVX1_RVT U557 ( .A(n491), .Y(n492) );
  INVX1_RVT U558 ( .A(\u_div/CryTmp[26][4] ), .Y(n491) );
  INVX1_RVT U559 ( .A(n541), .Y(n572) );
  INVX1_RVT U560 ( .A(n781), .Y(\u_div/PartRem[8][1] ) );
  INVX1_RVT U561 ( .A(\u_div/CryTmp[6][4] ), .Y(n877) );
  IBUFFX4_RVT U562 ( .A(n540), .Y(\u_div/PartRem[21][9] ) );
  INVX1_RVT U563 ( .A(net29601), .Y(\u_div/PartRem[9][6] ) );
  INVX1_RVT U564 ( .A(n879), .Y(n880) );
  INVX1_RVT U565 ( .A(n877), .Y(n878) );
  INVX1_RVT U566 ( .A(\u_div/PartRem[7][4] ), .Y(n879) );
  INVX1_RVT U567 ( .A(n881), .Y(n882) );
  INVX1_RVT U568 ( .A(\u_div/PartRem[7][5] ), .Y(n881) );
  INVX1_RVT U569 ( .A(net30407), .Y(\u_div/PartRem[10][8] ) );
  INVX1_RVT U570 ( .A(n784), .Y(\u_div/PartRem[7][3] ) );
  MUX21X1_RVT U571 ( .A1(net29676), .A2(net30288), .S0(quotient[5]), .Y(n856)
         );
  INVX1_RVT U572 ( .A(n848), .Y(n849) );
  INVX1_RVT U573 ( .A(\u_div/CryTmp[5][5] ), .Y(n848) );
  NAND2X0_RVT U574 ( .A1(net45599), .A2(\u_div/SumTmp[5][0] ), .Y(n1043) );
  INVX1_RVT U575 ( .A(net29674), .Y(\u_div/PartRem[6][6] ) );
  INVX1_RVT U576 ( .A(n852), .Y(n853) );
  INVX1_RVT U577 ( .A(\u_div/CryTmp[6][6] ), .Y(n852) );
  INVX1_RVT U578 ( .A(n850), .Y(n851) );
  INVX1_RVT U579 ( .A(\u_div/CryTmp[5][6] ), .Y(n850) );
  INVX1_RVT U580 ( .A(net51994), .Y(n787) );
  MUX21X1_RVT U581 ( .A1(\u_div/PartRem[7][6] ), .A2(\u_div/SumTmp[6][6] ), 
        .S0(net45257), .Y(net51994) );
  INVX1_RVT U582 ( .A(n509), .Y(n510) );
  INVX1_RVT U583 ( .A(\u_div/CryTmp[24][10] ), .Y(n509) );
  INVX1_RVT U584 ( .A(\u_div/SumTmp[26][9] ), .Y(net30830) );
  INVX1_RVT U585 ( .A(n520), .Y(n521) );
  INVX1_RVT U586 ( .A(\u_div/CryTmp[25][9] ), .Y(n520) );
  INVX1_RVT U587 ( .A(net40783), .Y(net29622) );
  INVX1_RVT U588 ( .A(\u_div/SumTmp[5][4] ), .Y(net30288) );
  INVX1_RVT U589 ( .A(n840), .Y(n841) );
  INVX1_RVT U590 ( .A(n856), .Y(\u_div/PartRem[5][5] ) );
  INVX1_RVT U591 ( .A(\u_div/CryTmp[4][5] ), .Y(n840) );
  INVX1_RVT U592 ( .A(\u_div/SumTmp[3][3] ), .Y(net30311) );
  INVX1_RVT U593 ( .A(\u_div/SumTmp[4][4] ), .Y(net30297) );
  INVX1_RVT U594 ( .A(\u_div/SumTmp[3][4] ), .Y(net30304) );
  INVX1_RVT U595 ( .A(n1036), .Y(\u_div/PartRem[3][5] ) );
  INVX1_RVT U596 ( .A(net49608), .Y(n804) );
  MUX21X1_RVT U597 ( .A1(\u_div/PartRem[6][6] ), .A2(\u_div/SumTmp[5][6] ), 
        .S0(net49616), .Y(net49608) );
  INVX1_RVT U598 ( .A(n804), .Y(n869) );
  INVX1_RVT U599 ( .A(\u_div/CryTmp[4][7] ), .Y(n866) );
  INVX1_RVT U600 ( .A(n842), .Y(net42516) );
  INVX2_RVT U601 ( .A(n455), .Y(n456) );
  IBUFFX4_RVT U602 ( .A(\u_div/SumTmp[13][12] ), .Y(net31123) );
  INVX0_RVT U603 ( .A(b[0]), .Y(net32406) );
  INVX2_RVT U604 ( .A(net49112), .Y(net49113) );
  INVX1_RVT U605 ( .A(net46962), .Y(net44969) );
  INVX0_RVT U606 ( .A(net32544), .Y(net49094) );
  INVX1_RVT U607 ( .A(\u_div/PartRem[11][11] ), .Y(n750) );
  INVX1_RVT U608 ( .A(n771), .Y(n772) );
  INVX1_RVT U609 ( .A(\u_div/CryTmp[8][10] ), .Y(n771) );
  INVX1_RVT U610 ( .A(net49280), .Y(net49281) );
  INVX1_RVT U611 ( .A(\u_div/CryTmp[6][10] ), .Y(net49280) );
  MUX21X1_RVT U612 ( .A1(\u_div/SumTmp[6][9] ), .A2(n876), .S0(net52013), .Y(
        n875) );
  INVX1_RVT U613 ( .A(n782), .Y(n876) );
  INVX1_RVT U614 ( .A(\u_div/CryTmp[3][10] ), .Y(n860) );
  MUX21X1_RVT U615 ( .A1(net29702), .A2(net30287), .S0(net42034), .Y(net29729)
         );
  INVX1_RVT U616 ( .A(\u_div/SumTmp[4][5] ), .Y(net30287) );
  MUX21X1_RVT U617 ( .A1(net29676), .A2(net30288), .S0(net44755), .Y(net29702)
         );
  INVX1_RVT U618 ( .A(net42516), .Y(net42520) );
  INVX1_RVT U619 ( .A(net29729), .Y(\u_div/PartRem[4][6] ) );
  INVX1_RVT U620 ( .A(\u_div/SumTmp[4][6] ), .Y(net30472) );
  INVX1_RVT U621 ( .A(n1033), .Y(\u_div/PartRem[3][8] ) );
  INVX1_RVT U622 ( .A(\u_div/CryTmp[2][8] ), .Y(n956) );
  INVX1_RVT U623 ( .A(n1035), .Y(\u_div/PartRem[3][6] ) );
  INVX1_RVT U624 ( .A(\u_div/CryTmp[2][6] ), .Y(n996) );
  NBUFFX2_RVT U625 ( .A(net42519), .Y(net45582) );
  INVX1_RVT U626 ( .A(net42516), .Y(net42519) );
  MUX21X1_RVT U627 ( .A1(n804), .A2(net30462), .S0(net50726), .Y(net29727) );
  INVX1_RVT U628 ( .A(\u_div/SumTmp[4][7] ), .Y(net30462) );
  INVX1_RVT U629 ( .A(n845), .Y(n846) );
  INVX1_RVT U630 ( .A(\u_div/CryTmp[3][8] ), .Y(n845) );
  INVX1_RVT U631 ( .A(net45228), .Y(net45229) );
  INVX1_RVT U632 ( .A(net30452), .Y(net45228) );
  INVX1_RVT U633 ( .A(\u_div/SumTmp[4][8] ), .Y(net30452) );
  INVX1_RVT U634 ( .A(net42516), .Y(net42517) );
  INVX1_RVT U635 ( .A(net30003), .Y(\u_div/PartRem[27][10] ) );
  INVX1_RVT U636 ( .A(\u_div/SumTmp[27][10] ), .Y(net30735) );
  INVX1_RVT U637 ( .A(net29983), .Y(\u_div/PartRem[28][10] ) );
  INVX1_RVT U638 ( .A(n875), .Y(n802) );
  INVX1_RVT U639 ( .A(net52003), .Y(net29671) );
  INVX1_RVT U640 ( .A(n860), .Y(n861) );
  INVX1_RVT U641 ( .A(n1034), .Y(\u_div/PartRem[3][7] ) );
  MUX21X1_RVT U642 ( .A1(net29729), .A2(net30286), .S0(net45584), .Y(n1034) );
  NBUFFX2_RVT U643 ( .A(net42520), .Y(net45581) );
  INVX1_RVT U644 ( .A(\u_div/SumTmp[3][6] ), .Y(net30286) );
  MUX21X1_RVT U645 ( .A1(net29728), .A2(net30471), .S0(net45585), .Y(n1033) );
  INVX1_RVT U646 ( .A(\u_div/SumTmp[3][7] ), .Y(net30471) );
  INVX1_RVT U647 ( .A(n935), .Y(n936) );
  INVX1_RVT U648 ( .A(n956), .Y(n957) );
  NBUFFX2_RVT U649 ( .A(net45582), .Y(net45583) );
  INVX1_RVT U650 ( .A(\u_div/SumTmp[3][8] ), .Y(net30461) );
  INVX1_RVT U651 ( .A(n1032), .Y(\u_div/PartRem[3][9] ) );
  INVX1_RVT U652 ( .A(net52000), .Y(net29672) );
  NBUFFX2_RVT U653 ( .A(net30442), .Y(net46608) );
  INVX1_RVT U654 ( .A(\u_div/SumTmp[4][9] ), .Y(net30442) );
  INVX1_RVT U655 ( .A(net42548), .Y(net42514) );
  INVX1_RVT U656 ( .A(\u_div/SumTmp[3][10] ), .Y(net30441) );
  INVX1_RVT U657 ( .A(n1053), .Y(\u_div/PartRem[3][10] ) );
  MUX21X1_RVT U658 ( .A1(net29726), .A2(net30451), .S0(net45587), .Y(n1053) );
  NBUFFX2_RVT U659 ( .A(net42517), .Y(net45584) );
  INVX1_RVT U660 ( .A(\u_div/SumTmp[3][9] ), .Y(net30451) );
  INVX2_RVT U661 ( .A(n513), .Y(n514) );
  INVX1_RVT U662 ( .A(n457), .Y(\u_div/PartRem[30][8] ) );
  NBUFFX2_RVT U663 ( .A(n569), .Y(n575) );
  INVX2_RVT U664 ( .A(n162), .Y(n630) );
  INVX1_RVT U665 ( .A(n493), .Y(n495) );
  INVX1_RVT U666 ( .A(\u_div/CryTmp[26][11] ), .Y(n493) );
  INVX1_RVT U667 ( .A(n1003), .Y(n1026) );
  INVX1_RVT U668 ( .A(net29752), .Y(\u_div/PartRem[4][12] ) );
  MUX21X1_RVT U669 ( .A1(\u_div/PartRem[3][7] ), .A2(\u_div/SumTmp[2][7] ), 
        .S0(n987), .Y(n951) );
  INVX1_RVT U670 ( .A(n998), .Y(n999) );
  INVX1_RVT U671 ( .A(\u_div/CryTmp[1][8] ), .Y(n998) );
  INVX1_RVT U672 ( .A(n1174), .Y(\u_div/PartRem[2][9] ) );
  INVX1_RVT U673 ( .A(\u_div/CryTmp[1][9] ), .Y(n954) );
  MUX21X1_RVT U674 ( .A1(n1032), .A2(n1173), .S0(n953), .Y(n1172) );
  INVX1_RVT U675 ( .A(n1052), .Y(n1011) );
  NBUFFX2_RVT U676 ( .A(net42514), .Y(net45585) );
  MUX21X1_RVT U677 ( .A1(\u_div/PartRem[3][10] ), .A2(\u_div/SumTmp[2][10] ), 
        .S0(quotient[2]), .Y(n982) );
  INVX1_RVT U678 ( .A(net30063), .Y(\u_div/PartRem[24][15] ) );
  IBUFFX4_RVT U679 ( .A(n1098), .Y(\u_div/PartRem[23][15] ) );
  MUX21X1_RVT U680 ( .A1(net30041), .A2(net30636), .S0(net47709), .Y(n532) );
  INVX1_RVT U681 ( .A(n532), .Y(\u_div/PartRem[24][16] ) );
  MUX21X1_RVT U682 ( .A1(net49255), .A2(net30356), .S0(net40719), .Y(n1022) );
  INVX1_RVT U683 ( .A(net29751), .Y(\u_div/PartRem[4][13] ) );
  INVX1_RVT U684 ( .A(\u_div/CryTmp[1][14] ), .Y(n915) );
  INVX1_RVT U685 ( .A(net29820), .Y(\u_div/PartRem[39][1] ) );
  INVX1_RVT U686 ( .A(n566), .Y(n573) );
  INVX1_RVT U687 ( .A(\u_div/CryTmp[23][17] ), .Y(n566) );
  INVX1_RVT U688 ( .A(\u_div/CryTmp[10][16] ), .Y(n303) );
  INVX1_RVT U689 ( .A(n964), .Y(n1058) );
  INVX0_RVT U690 ( .A(net29980), .Y(\u_div/PartRem[28][13] ) );
  INVX1_RVT U691 ( .A(n864), .Y(n865) );
  INVX1_RVT U692 ( .A(\u_div/CryTmp[3][14] ), .Y(n864) );
  INVX1_RVT U693 ( .A(n1048), .Y(\u_div/PartRem[3][15] ) );
  INVX1_RVT U694 ( .A(n1168), .Y(\u_div/PartRem[2][14] ) );
  MUX21X1_RVT U695 ( .A1(n1050), .A2(n1169), .S0(n953), .Y(n1168) );
  INVX1_RVT U696 ( .A(\u_div/SumTmp[2][13] ), .Y(n1169) );
  INVX1_RVT U697 ( .A(n923), .Y(n924) );
  IBUFFX4_RVT U698 ( .A(n916), .Y(n923) );
  INVX1_RVT U699 ( .A(\u_div/CryTmp[1][13] ), .Y(n913) );
  INVX0_RVT U700 ( .A(n1058), .Y(n888) );
  IBUFFX4_RVT U701 ( .A(net30123), .Y(\u_div/PartRem[23][17] ) );
  INVX1_RVT U702 ( .A(n574), .Y(n567) );
  INVX1_RVT U703 ( .A(n573), .Y(n574) );
  MUX21X1_RVT U704 ( .A1(net30039), .A2(net30540), .S0(net47709), .Y(n530) );
  INVX1_RVT U705 ( .A(n609), .Y(n633) );
  MUX21X1_RVT U706 ( .A1(net30659), .A2(net30977), .S0(n45), .Y(n691) );
  MUX21X1_RVT U707 ( .A1(net29664), .A2(net30354), .S0(net40656), .Y(n795) );
  INVX1_RVT U708 ( .A(net42548), .Y(net42515) );
  INVX1_RVT U709 ( .A(n919), .Y(n903) );
  INVX1_RVT U710 ( .A(\u_div/CryTmp[2][16] ), .Y(n919) );
  INVX1_RVT U711 ( .A(n971), .Y(n972) );
  INVX1_RVT U712 ( .A(\u_div/CryTmp[0][15] ), .Y(n976) );
  INVX1_RVT U713 ( .A(net29782), .Y(\u_div/PartRem[40][1] ) );
  IBUFFX4_RVT U714 ( .A(net30181), .Y(\u_div/PartRem[22][18] ) );
  XOR2X1_RVT U715 ( .A1(\u_div/PartRem[8][18] ), .A2(net31940), .Y(n1002) );
  INVX1_RVT U716 ( .A(n858), .Y(n871) );
  INVX1_RVT U717 ( .A(\u_div/CryTmp[4][21] ), .Y(n858) );
  INVX0_RVT U718 ( .A(net40656), .Y(net45737) );
  INVX1_RVT U719 ( .A(\u_div/PartRem[38][4] ), .Y(n988) );
  MUX21X1_RVT U720 ( .A1(\u_div/SumTmp[5][21] ), .A2(\u_div/PartRem[6][21] ), 
        .S0(net45654), .Y(n873) );
  INVX2_RVT U721 ( .A(n884), .Y(n885) );
  INVX1_RVT U722 ( .A(n904), .Y(n920) );
  INVX1_RVT U723 ( .A(n903), .Y(n904) );
  IBUFFX4_RVT U724 ( .A(\u_div/PartRem[1][17] ), .Y(n965) );
  INVX1_RVT U725 ( .A(n969), .Y(n970) );
  INVX1_RVT U726 ( .A(\u_div/PartRem[33][11] ), .Y(n325) );
  IBUFFX4_RVT U727 ( .A(\u_div/SumTmp[34][8] ), .Y(n429) );
  INVX1_RVT U728 ( .A(\u_div/PartRem[35][8] ), .Y(net46238) );
  IBUFFX4_RVT U729 ( .A(net29818), .Y(\u_div/PartRem[39][3] ) );
  MUX21X1_RVT U730 ( .A1(net30799), .A2(net31021), .S0(net32548), .Y(net30845)
         );
  MUX21X1_RVT U731 ( .A1(n791), .A2(n824), .S0(quotient[5]), .Y(n809) );
  INVX1_RVT U732 ( .A(\u_div/SumTmp[5][20] ), .Y(n824) );
  INVX1_RVT U733 ( .A(n872), .Y(n859) );
  INVX1_RVT U734 ( .A(n809), .Y(\u_div/PartRem[5][21] ) );
  INVX1_RVT U735 ( .A(n871), .Y(n872) );
  INVX1_RVT U736 ( .A(net29684), .Y(net38272) );
  INVX1_RVT U737 ( .A(net52012), .Y(net52013) );
  INVX1_RVT U738 ( .A(net45737), .Y(net52012) );
  INVX2_RVT U739 ( .A(n238), .Y(n632) );
  INVX1_RVT U740 ( .A(net30657), .Y(\u_div/PartRem[16][19] ) );
  INVX1_RVT U741 ( .A(net50742), .Y(net50743) );
  INVX1_RVT U742 ( .A(net38274), .Y(net50742) );
  INVX1_RVT U743 ( .A(n793), .Y(\u_div/PartRem[6][19] ) );
  NBUFFX2_RVT U744 ( .A(\u_div/PartRem[4][19] ), .Y(n857) );
  INVX1_RVT U745 ( .A(n822), .Y(\u_div/PartRem[4][19] ) );
  INVX1_RVT U746 ( .A(n945), .Y(n946) );
  INVX1_RVT U747 ( .A(\u_div/CryTmp[0][18] ), .Y(n945) );
  NBUFFX2_RVT U748 ( .A(net42523), .Y(net45592) );
  INVX1_RVT U749 ( .A(net42548), .Y(net42523) );
  INVX2_RVT U750 ( .A(n442), .Y(n449) );
  INVX1_RVT U751 ( .A(\u_div/PartRem[31][13] ), .Y(n451) );
  INVX1_RVT U752 ( .A(\u_div/CryTmp[31][13] ), .Y(n440) );
  INVX1_RVT U753 ( .A(n325), .Y(n326) );
  INVX1_RVT U754 ( .A(n963), .Y(n1055) );
  MUX21X1_RVT U755 ( .A1(\u_div/SumTmp[38][5] ), .A2(\u_div/PartRem[39][5] ), 
        .S0(net46142), .Y(n963) );
  INVX1_RVT U756 ( .A(net29741), .Y(\u_div/PartRem[4][22] ) );
  MUX21X1_RVT U757 ( .A1(net38272), .A2(\u_div/SumTmp[5][22] ), .S0(net44755), 
        .Y(n836) );
  INVX1_RVT U758 ( .A(n311), .Y(n312) );
  INVX1_RVT U759 ( .A(net52013), .Y(net45257) );
  MUX21X1_RVT U760 ( .A1(net50743), .A2(\u_div/SumTmp[3][23] ), .S0(net45583), 
        .Y(\u_div/PartRem[3][24] ) );
  INVX1_RVT U761 ( .A(net30016), .Y(\u_div/PartRem[26][18] ) );
  NBUFFX2_RVT U762 ( .A(\u_div/CryTmp[4][20] ), .Y(n870) );
  INVX1_RVT U763 ( .A(n941), .Y(n942) );
  INVX1_RVT U764 ( .A(\u_div/CryTmp[0][19] ), .Y(n941) );
  INVX1_RVT U765 ( .A(n450), .Y(n443) );
  INVX2_RVT U766 ( .A(n451), .Y(n452) );
  INVX1_RVT U767 ( .A(net29815), .Y(\u_div/PartRem[39][6] ) );
  INVX1_RVT U768 ( .A(n962), .Y(n1054) );
  MUX21X1_RVT U769 ( .A1(\u_div/PartRem[39][6] ), .A2(\u_div/SumTmp[38][6] ), 
        .S0(net37581), .Y(n962) );
  IBUFFX4_RVT U770 ( .A(net30177), .Y(\u_div/PartRem[22][21] ) );
  IBUFFX4_RVT U771 ( .A(n1120), .Y(\u_div/PartRem[22][23] ) );
  INVX1_RVT U772 ( .A(net30117), .Y(\u_div/PartRem[23][22] ) );
  IBUFFX4_RVT U773 ( .A(n526), .Y(\u_div/PartRem[24][21] ) );
  INVX1_RVT U774 ( .A(\u_div/SumTmp[8][21] ), .Y(net29681) );
  INVX1_RVT U775 ( .A(n1072), .Y(\u_div/PartRem[3][23] ) );
  INVX1_RVT U776 ( .A(\u_div/SumTmp[3][22] ), .Y(net29939) );
  NOR2X1_RVT U777 ( .A1(\u_div/CryTmp[3][24] ), .A2(\u_div/PartRem[4][24] ), 
        .Y(net45183) );
  MUX21X1_RVT U778 ( .A1(\u_div/SumTmp[4][23] ), .A2(n836), .S0(net38350), .Y(
        \u_div/PartRem[4][24] ) );
  INVX1_RVT U779 ( .A(n980), .Y(n981) );
  INVX1_RVT U780 ( .A(n985), .Y(n980) );
  INVX1_RVT U781 ( .A(n1008), .Y(n1015) );
  INVX1_RVT U782 ( .A(\u_div/SumTmp[27][17] ), .Y(net30204) );
  INVX1_RVT U783 ( .A(n890), .Y(n987) );
  INVX1_RVT U784 ( .A(\u_div/CryTmp[0][21] ), .Y(n925) );
  MUX21X1_RVT U785 ( .A1(n1019), .A2(n1020), .S0(net32530), .Y(net29628) );
  MUX21X1_RVT U786 ( .A1(net30118), .A2(net30247), .S0(net32610), .Y(n1119) );
  INVX1_RVT U787 ( .A(net38343), .Y(net32596) );
  IBUFFX4_RVT U788 ( .A(net51611), .Y(net51612) );
  INVX1_RVT U789 ( .A(n1019), .Y(\u_div/PartRem[10][22] ) );
  INVX1_RVT U790 ( .A(\u_div/PartRem[38][8] ), .Y(net44464) );
  INVX2_RVT U791 ( .A(net42357), .Y(net32560) );
  INVX1_RVT U792 ( .A(net30653), .Y(\u_div/PartRem[16][22] ) );
  MUX21X1_RVT U793 ( .A1(\u_div/PartRem[19][22] ), .A2(\u_div/SumTmp[18][22] ), 
        .S0(net45671), .Y(n638) );
  MUX21X1_RVT U794 ( .A1(net29975), .A2(net30144), .S0(net41415), .Y(net29994)
         );
  INVX1_RVT U795 ( .A(\u_div/SumTmp[3][21] ), .Y(net30331) );
  INVX1_RVT U796 ( .A(n1041), .Y(\u_div/PartRem[3][22] ) );
  INVX1_RVT U797 ( .A(n987), .Y(n952) );
  INVX1_RVT U798 ( .A(n912), .Y(n979) );
  INVX1_RVT U799 ( .A(n911), .Y(n912) );
  INVX1_RVT U800 ( .A(n978), .Y(n911) );
  IBUFFX4_RVT U801 ( .A(\u_div/CryTmp[1][23] ), .Y(n978) );
  INVX1_RVT U802 ( .A(\u_div/CryTmp[0][22] ), .Y(n921) );
  INVX1_RVT U803 ( .A(n925), .Y(n926) );
  IBUFFX4_RVT U804 ( .A(\u_div/CryTmp[24][22] ), .Y(net48533) );
  IBUFFX16_RVT U805 ( .A(n423), .Y(\u_div/PartRem[31][15] ) );
  INVX1_RVT U806 ( .A(net31297), .Y(net39870) );
  INVX1_RVT U807 ( .A(n350), .Y(\u_div/PartRem[39][8] ) );
  INVX1_RVT U808 ( .A(net42040), .Y(net42041) );
  INVX1_RVT U809 ( .A(n967), .Y(n968) );
  NBUFFX8_RVT U810 ( .A(net32130), .Y(net49055) );
  INVX1_RVT U811 ( .A(net30675), .Y(\u_div/PartRem[16][23] ) );
  INVX2_RVT U812 ( .A(n293), .Y(n294) );
  IBUFFX4_RVT U813 ( .A(\u_div/PartRem[1][23] ), .Y(n907) );
  MUX21X1_RVT U814 ( .A1(n1041), .A2(n1143), .S0(n953), .Y(n1142) );
  INVX0_RVT U815 ( .A(net31814), .Y(net31800) );
  INVX1_RVT U816 ( .A(n921), .Y(n922) );
  IBUFFX4_RVT U817 ( .A(\u_div/PartRem[1][22] ), .Y(n909) );
  INVX1_RVT U818 ( .A(net52992), .Y(net48534) );
  INVX0_RVT U819 ( .A(net32024), .Y(net52311) );
  INVX1_RVT U820 ( .A(net45007), .Y(net32598) );
  INVX2_RVT U821 ( .A(n560), .Y(net32610) );
  INVX1_RVT U822 ( .A(net42041), .Y(net42034) );
  INVX1_RVT U823 ( .A(net45669), .Y(net45665) );
  INVX1_RVT U824 ( .A(n232), .Y(net48658) );
  IBUFFX4_RVT U825 ( .A(net44394), .Y(net44395) );
  INVX1_RVT U826 ( .A(net29992), .Y(\u_div/PartRem[27][20] ) );
  MUX21X1_RVT U827 ( .A1(\u_div/PartRem[2][23] ), .A2(\u_div/SumTmp[1][23] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][24] ) );
  NOR2X1_RVT U828 ( .A1(net31287), .A2(net31291), .Y(net37563) );
  IBUFFX4_RVT U829 ( .A(\u_div/CryTmp[34][13] ), .Y(net31291) );
  NBUFFX4_RVT U830 ( .A(net37556), .Y(net43819) );
  INVX1_RVT U831 ( .A(net48658), .Y(net48659) );
  AND2X1_RVT U832 ( .A1(n1006), .A2(\u_div/CryTmp[35][12] ), .Y(net37585) );
  INVX1_RVT U833 ( .A(\u_div/CryTmp[36][11] ), .Y(net31281) );
  INVX2_RVT U834 ( .A(n375), .Y(n376) );
  IBUFFX4_RVT U835 ( .A(net30069), .Y(\u_div/PartRem[23][9] ) );
  MUX21X2_RVT U836 ( .A1(net30188), .A2(net30983), .S0(n191), .Y(n553) );
  IBUFFX4_RVT U837 ( .A(net30070), .Y(\u_div/PartRem[23][8] ) );
  INVX2_RVT U838 ( .A(n242), .Y(n564) );
  IBUFFX16_RVT U839 ( .A(net30283), .Y(\u_div/PartRem[20][10] ) );
  IBUFFX2_RVT U840 ( .A(n551), .Y(\u_div/PartRem[21][14] ) );
  INVX2_RVT U841 ( .A(n556), .Y(\u_div/PartRem[20][17] ) );
  AND3X2_RVT U842 ( .A1(\u_div/CryTmp[39][8] ), .A2(net32198), .A3(net37169), 
        .Y(net47716) );
  MUX21X2_RVT U843 ( .A1(n418), .A2(n425), .S0(net50049), .Y(net29900) );
  INVX32_RVT U844 ( .A(net30002), .Y(n281) );
  IBUFFX16_RVT U845 ( .A(n281), .Y(n282) );
  INVX2_RVT U846 ( .A(n282), .Y(\u_div/PartRem[27][11] ) );
  MUX21X2_RVT U847 ( .A1(n282), .A2(net30734), .S0(n152), .Y(net30022) );
  IBUFFX16_RVT U848 ( .A(\u_div/SumTmp[31][5] ), .Y(net30787) );
  IBUFFX4_RVT U849 ( .A(\u_div/CryTmp[31][8] ), .Y(n436) );
  INVX1_RVT U850 ( .A(\u_div/SumTmp[37][2] ), .Y(n362) );
  MUX21X2_RVT U851 ( .A1(net30846), .A2(net31042), .S0(net32544), .Y(net30892)
         );
  IBUFFX4_RVT U852 ( .A(\u_div/SumTmp[11][18] ), .Y(net31042) );
  IBUFFX4_RVT U853 ( .A(net30890), .Y(\u_div/PartRem[11][20] ) );
  INVX4_RVT U854 ( .A(n649), .Y(\u_div/PartRem[17][5] ) );
  MUX21X2_RVT U855 ( .A1(net30531), .A2(net31188), .S0(net32580), .Y(n649) );
  MUX21X2_RVT U856 ( .A1(net45288), .A2(net31064), .S0(net32542), .Y(net30893)
         );
  MUX21X2_RVT U857 ( .A1(net30842), .A2(net30973), .S0(net32542), .Y(net30888)
         );
  INVX1_RVT U858 ( .A(net38336), .Y(net32542) );
  OR2X2_RVT U859 ( .A1(\u_div/PartRem[19][24] ), .A2(\u_div/CryTmp[18][24] ), 
        .Y(n635) );
  INVX4_RVT U860 ( .A(n634), .Y(net45669) );
  OR2X2_RVT U861 ( .A1(\u_div/PartRem[19][24] ), .A2(\u_div/CryTmp[18][24] ), 
        .Y(n634) );
  IBUFFX2_RVT U862 ( .A(\u_div/CryTmp[36][9] ), .Y(n283) );
  IBUFFX4_RVT U863 ( .A(n283), .Y(n284) );
  INVX8_RVT U864 ( .A(b[9]), .Y(net32186) );
  MUX21X1_RVT U865 ( .A1(n1065), .A2(n1084), .S0(net37570), .Y(n1068) );
  IBUFFX16_RVT U866 ( .A(\u_div/SumTmp[37][6] ), .Y(n1128) );
  IBUFFX16_RVT U867 ( .A(n1065), .Y(\u_div/PartRem[37][10] ) );
  IBUFFX4_RVT U868 ( .A(n394), .Y(\u_div/PartRem[35][5] ) );
  INVX2_RVT U869 ( .A(net31107), .Y(n285) );
  INVX1_RVT U870 ( .A(n285), .Y(n286) );
  IBUFFX16_RVT U871 ( .A(\u_div/CryTmp[16][5] ), .Y(n287) );
  INVX4_RVT U872 ( .A(n287), .Y(n288) );
  IBUFFX4_RVT U873 ( .A(net30071), .Y(\u_div/PartRem[23][7] ) );
  IBUFFX4_RVT U874 ( .A(net30072), .Y(\u_div/PartRem[23][6] ) );
  IBUFFX4_RVT U875 ( .A(n533), .Y(\u_div/PartRem[23][5] ) );
  IBUFFX4_RVT U876 ( .A(n534), .Y(\u_div/PartRem[23][3] ) );
  IBUFFX4_RVT U877 ( .A(n535), .Y(\u_div/PartRem[23][2] ) );
  IBUFFX16_RVT U878 ( .A(\u_div/CryTmp[25][19] ), .Y(n291) );
  IBUFFX16_RVT U879 ( .A(\u_div/CryTmp[25][21] ), .Y(n293) );
  IBUFFX16_RVT U880 ( .A(\u_div/CryTmp[17][22] ), .Y(n295) );
  INVX4_RVT U881 ( .A(n295), .Y(n296) );
  IBUFFX16_RVT U882 ( .A(net30664), .Y(\u_div/PartRem[16][12] ) );
  IBUFFX4_RVT U883 ( .A(net30663), .Y(\u_div/PartRem[16][13] ) );
  MUX21X1_RVT U884 ( .A1(net30665), .A2(n286), .S0(n58), .Y(n663) );
  INVX4_RVT U885 ( .A(n746), .Y(n747) );
  IBUFFX16_RVT U886 ( .A(\u_div/CryTmp[15][12] ), .Y(n297) );
  INVX4_RVT U887 ( .A(n297), .Y(n298) );
  IBUFFX4_RVT U888 ( .A(\u_div/SumTmp[16][14] ), .Y(net31025) );
  IBUFFX4_RVT U889 ( .A(net30021), .Y(\u_div/PartRem[26][13] ) );
  IBUFFX4_RVT U890 ( .A(net30662), .Y(\u_div/PartRem[16][14] ) );
  IBUFFX16_RVT U891 ( .A(\u_div/CryTmp[10][20] ), .Y(n299) );
  INVX4_RVT U892 ( .A(n299), .Y(n300) );
  IBUFFX16_RVT U893 ( .A(\u_div/CryTmp[9][11] ), .Y(n301) );
  INVX4_RVT U894 ( .A(n301), .Y(n302) );
  IBUFFX4_RVT U895 ( .A(n303), .Y(n304) );
  IBUFFX16_RVT U896 ( .A(net30895), .Y(\u_div/PartRem[11][16] ) );
  INVX2_RVT U897 ( .A(n349), .Y(\u_div/PartRem[40][2] ) );
  IBUFFX16_RVT U898 ( .A(\u_div/CryTmp[43][2] ), .Y(n307) );
  INVX4_RVT U899 ( .A(n307), .Y(n308) );
  IBUFFX4_RVT U900 ( .A(n552), .Y(\u_div/PartRem[21][13] ) );
  IBUFFX16_RVT U901 ( .A(net30187), .Y(\u_div/PartRem[22][12] ) );
  INVX4_RVT U902 ( .A(n568), .Y(n569) );
  IBUFFX16_RVT U903 ( .A(net30131), .Y(\u_div/PartRem[22][9] ) );
  IBUFFX16_RVT U904 ( .A(n553), .Y(\u_div/PartRem[21][12] ) );
  IBUFFX4_RVT U905 ( .A(n593), .Y(\u_div/PartRem[21][19] ) );
  INVX32_RVT U906 ( .A(\u_div/CryTmp[20][11] ), .Y(n309) );
  IBUFFX16_RVT U907 ( .A(n309), .Y(n310) );
  IBUFFX16_RVT U908 ( .A(n554), .Y(\u_div/PartRem[21][11] ) );
  MUX21X2_RVT U909 ( .A1(net30132), .A2(net31052), .S0(n205), .Y(n540) );
  INVX8_RVT U910 ( .A(b[7]), .Y(net32242) );
  IBUFFX16_RVT U911 ( .A(net30132), .Y(\u_div/PartRem[22][8] ) );
  IBUFFX4_RVT U912 ( .A(net29934), .Y(\u_div/PartRem[30][13] ) );
  IBUFFX4_RVT U913 ( .A(\u_div/CryTmp[26][21] ), .Y(n484) );
  IBUFFX4_RVT U914 ( .A(\u_div/CryTmp[11][20] ), .Y(n311) );
  INVX2_RVT U915 ( .A(n692), .Y(\u_div/PartRem[15][17] ) );
  IBUFFX16_RVT U916 ( .A(\u_div/CryTmp[14][16] ), .Y(n746) );
  INVX0_RVT U917 ( .A(n693), .Y(\u_div/PartRem[15][16] ) );
  MUX21X1_RVT U918 ( .A1(net30133), .A2(net31074), .S0(n201), .Y(n541) );
  IBUFFX16_RVT U919 ( .A(\u_div/SumTmp[7][20] ), .Y(net29737) );
  IBUFFX32_RVT U920 ( .A(n1028), .Y(\u_div/PartRem[7][22] ) );
  XOR3X1_RVT U921 ( .A1(\u_div/PartRem[2][23] ), .A2(n979), .A3(net31800), .Y(
        \u_div/SumTmp[1][23] ) );
  IBUFFX16_RVT U922 ( .A(net30133), .Y(\u_div/PartRem[22][7] ) );
  IBUFFX16_RVT U923 ( .A(\u_div/CryTmp[21][7] ), .Y(n313) );
  INVX4_RVT U924 ( .A(n313), .Y(n314) );
  IBUFFX16_RVT U925 ( .A(net30417), .Y(\u_div/PartRem[10][7] ) );
  IBUFFX16_RVT U926 ( .A(\u_div/CryTmp[9][7] ), .Y(n315) );
  INVX4_RVT U927 ( .A(n315), .Y(n316) );
  IBUFFX16_RVT U928 ( .A(\u_div/CryTmp[15][21] ), .Y(n317) );
  IBUFFX16_RVT U929 ( .A(\u_div/CryTmp[15][20] ), .Y(n319) );
  INVX4_RVT U930 ( .A(n319), .Y(n320) );
  INVX1_RVT U931 ( .A(n518), .Y(n519) );
  IBUFFX4_RVT U932 ( .A(\u_div/CryTmp[25][13] ), .Y(n518) );
  IBUFFX16_RVT U933 ( .A(\u_div/CryTmp[25][11] ), .Y(n321) );
  INVX4_RVT U934 ( .A(n321), .Y(n322) );
  INVX16_RVT U935 ( .A(\u_div/PartRem[28][17] ), .Y(n323) );
  IBUFFX4_RVT U936 ( .A(n323), .Y(n324) );
  INVX2_RVT U937 ( .A(n351), .Y(\u_div/PartRem[39][7] ) );
  INVX16_RVT U938 ( .A(net29633), .Y(\u_div/PartRem[8][20] ) );
  MUX21X1_RVT U939 ( .A1(\u_div/SumTmp[38][1] ), .A2(\u_div/PartRem[39][1] ), 
        .S0(net46142), .Y(net46015) );
  INVX1_RVT U940 ( .A(b[2]), .Y(net32368) );
  INVX1_RVT U941 ( .A(n352), .Y(\u_div/PartRem[38][1] ) );
  MUX21X1_RVT U942 ( .A1(net31546), .A2(net37262), .S0(net37581), .Y(n352) );
  INVX1_RVT U943 ( .A(b[1]), .Y(net32382) );
  OR2X1_RVT U944 ( .A1(net32408), .A2(a[37]), .Y(\u_div/CryTmp[37][1] ) );
  INVX8_RVT U945 ( .A(b[0]), .Y(net32408) );
  MUX21X1_RVT U946 ( .A1(net29828), .A2(n362), .S0(net37242), .Y(net29836) );
  IBUFFX16_RVT U947 ( .A(\u_div/CryTmp[37][3] ), .Y(net46241) );
  INVX0_RVT U948 ( .A(\u_div/SumTmp[37][1] ), .Y(net30697) );
  INVX1_RVT U949 ( .A(a[38]), .Y(net31546) );
  XOR2X1_RVT U950 ( .A1(a[38]), .A2(net32408), .Y(net37262) );
  AND2X1_RVT U951 ( .A1(net37169), .A2(\u_div/CryTmp[38][9] ), .Y(net37581) );
  MUX21X1_RVT U952 ( .A1(n352), .A2(net30697), .S0(net37242), .Y(net29837) );
  AND4X1_RVT U953 ( .A1(net31270), .A2(net31271), .A3(net31272), .A4(net31273), 
        .Y(net37169) );
  INVX1_RVT U954 ( .A(b[8]), .Y(net32212) );
  MUX21X1_RVT U955 ( .A1(n347), .A2(n359), .S0(quotient[39]), .Y(n351) );
  INVX2_RVT U956 ( .A(n381), .Y(n382) );
  IBUFFX16_RVT U957 ( .A(\u_div/CryTmp[38][7] ), .Y(n381) );
  INVX1_RVT U958 ( .A(b[6]), .Y(net32272) );
  INVX1_RVT U959 ( .A(net29816), .Y(\u_div/PartRem[39][5] ) );
  INVX1_RVT U960 ( .A(b[5]), .Y(net32302) );
  IBUFFX16_RVT U961 ( .A(net29817), .Y(\u_div/PartRem[39][4] ) );
  MUX21X1_RVT U962 ( .A1(n348), .A2(net30507), .S0(n171), .Y(net29817) );
  INVX1_RVT U963 ( .A(b[4]), .Y(net32326) );
  INVX32_RVT U964 ( .A(\u_div/CryTmp[38][4] ), .Y(n378) );
  MUX21X1_RVT U965 ( .A1(n349), .A2(net30555), .S0(n172), .Y(net29818) );
  OR2X1_RVT U966 ( .A1(net32408), .A2(a[38]), .Y(\u_div/CryTmp[38][1] ) );
  MUX21X1_RVT U967 ( .A1(\u_div/PartRem[39][8] ), .A2(\u_div/SumTmp[38][8] ), 
        .S0(net37581), .Y(net50339) );
  INVX0_RVT U968 ( .A(\u_div/SumTmp[38][7] ), .Y(n358) );
  MUX21X1_RVT U969 ( .A1(n341), .A2(net30157), .S0(net50182), .Y(n347) );
  INVX0_RVT U970 ( .A(\u_div/SumTmp[39][6] ), .Y(n359) );
  INVX1_RVT U971 ( .A(n347), .Y(\u_div/PartRem[40][6] ) );
  INVX1_RVT U972 ( .A(net29778), .Y(\u_div/PartRem[40][5] ) );
  MUX21X1_RVT U973 ( .A1(n342), .A2(net30217), .S0(net50182), .Y(net29778) );
  INVX1_RVT U974 ( .A(net29779), .Y(\u_div/PartRem[40][4] ) );
  MUX21X1_RVT U975 ( .A1(n343), .A2(net30265), .S0(n385), .Y(net29779) );
  INVX1_RVT U976 ( .A(n348), .Y(\u_div/PartRem[40][3] ) );
  MUX21X1_RVT U977 ( .A1(n344), .A2(net30508), .S0(net50186), .Y(n348) );
  INVX2_RVT U978 ( .A(n379), .Y(n380) );
  IBUFFX16_RVT U979 ( .A(\u_div/CryTmp[39][2] ), .Y(n379) );
  MUX21X1_RVT U980 ( .A1(net31514), .A2(net37252), .S0(net50182), .Y(net29782)
         );
  OR2X1_RVT U981 ( .A1(net32408), .A2(a[39]), .Y(\u_div/CryTmp[39][1] ) );
  MUX21X1_RVT U982 ( .A1(n351), .A2(n358), .S0(net37581), .Y(net29822) );
  INVX1_RVT U983 ( .A(n346), .Y(\u_div/PartRem[40][7] ) );
  MUX21X1_RVT U984 ( .A1(n340), .A2(n354), .S0(n385), .Y(n346) );
  INVX1_RVT U985 ( .A(net32210), .Y(net32198) );
  INVX0_RVT U986 ( .A(\u_div/SumTmp[39][7] ), .Y(n353) );
  MUX21X1_RVT U987 ( .A1(n336), .A2(n355), .S0(net37584), .Y(n340) );
  INVX0_RVT U988 ( .A(\u_div/SumTmp[40][6] ), .Y(n354) );
  IBUFFX4_RVT U989 ( .A(n340), .Y(\u_div/PartRem[41][6] ) );
  INVX1_RVT U990 ( .A(n341), .Y(\u_div/PartRem[41][5] ) );
  MUX21X1_RVT U991 ( .A1(n337), .A2(net30158), .S0(net37584), .Y(n341) );
  INVX1_RVT U992 ( .A(n342), .Y(\u_div/PartRem[41][4] ) );
  MUX21X1_RVT U993 ( .A1(n387), .A2(net30218), .S0(net37584), .Y(n342) );
  INVX1_RVT U994 ( .A(n343), .Y(\u_div/PartRem[41][3] ) );
  MUX21X1_RVT U995 ( .A1(n338), .A2(net30266), .S0(net37584), .Y(n343) );
  INVX1_RVT U996 ( .A(n344), .Y(\u_div/PartRem[41][2] ) );
  MUX21X1_RVT U997 ( .A1(n339), .A2(net30509), .S0(net37584), .Y(n344) );
  INVX2_RVT U998 ( .A(n345), .Y(\u_div/PartRem[41][1] ) );
  MUX21X1_RVT U999 ( .A1(net31498), .A2(net37256), .S0(net37584), .Y(n345) );
  OR2X1_RVT U1000 ( .A1(net32408), .A2(a[40]), .Y(\u_div/CryTmp[40][1] ) );
  MUX21X1_RVT U1001 ( .A1(n346), .A2(n353), .S0(n171), .Y(n350) );
  MUX21X1_RVT U1002 ( .A1(n332), .A2(n356), .S0(net43819), .Y(n336) );
  IBUFFX4_RVT U1003 ( .A(n336), .Y(\u_div/PartRem[42][5] ) );
  IBUFFX4_RVT U1004 ( .A(n337), .Y(\u_div/PartRem[42][4] ) );
  MUX21X1_RVT U1005 ( .A1(n333), .A2(net30159), .S0(net43819), .Y(n337) );
  IBUFFX4_RVT U1006 ( .A(n387), .Y(\u_div/PartRem[42][3] ) );
  IBUFFX16_RVT U1007 ( .A(n338), .Y(\u_div/PartRem[42][2] ) );
  INVX4_RVT U1008 ( .A(n383), .Y(n384) );
  IBUFFX16_RVT U1009 ( .A(\u_div/CryTmp[41][2] ), .Y(n383) );
  INVX2_RVT U1010 ( .A(n339), .Y(n377) );
  MUX21X2_RVT U1011 ( .A1(net31482), .A2(net37184), .S0(net37556), .Y(n339) );
  OR2X1_RVT U1012 ( .A1(net32408), .A2(a[41]), .Y(\u_div/CryTmp[41][1] ) );
  NOR2X4_RVT U1013 ( .A1(net31255), .A2(net43885), .Y(net37584) );
  MUX21X1_RVT U1014 ( .A1(n329), .A2(n357), .S0(quotient[43]), .Y(n332) );
  INVX0_RVT U1015 ( .A(\u_div/SumTmp[42][4] ), .Y(n356) );
  IBUFFX4_RVT U1016 ( .A(n333), .Y(\u_div/PartRem[43][3] ) );
  MUX21X1_RVT U1017 ( .A1(n330), .A2(n360), .S0(quotient[43]), .Y(n333) );
  MUX21X1_RVT U1018 ( .A1(n331), .A2(n361), .S0(quotient[43]), .Y(n334) );
  OR2X1_RVT U1019 ( .A1(net32408), .A2(a[42]), .Y(\u_div/CryTmp[42][1] ) );
  MUX21X1_RVT U1020 ( .A1(n327), .A2(net30098), .S0(quotient[44]), .Y(n329) );
  INVX1_RVT U1021 ( .A(n329), .Y(\u_div/PartRem[44][3] ) );
  IBUFFX16_RVT U1022 ( .A(n330), .Y(\u_div/PartRem[44][2] ) );
  MUX21X1_RVT U1023 ( .A1(n328), .A2(net30161), .S0(quotient[44]), .Y(n330) );
  INVX1_RVT U1024 ( .A(n331), .Y(\u_div/PartRem[44][1] ) );
  OR2X1_RVT U1025 ( .A1(net32408), .A2(a[43]), .Y(\u_div/CryTmp[43][1] ) );
  NOR3X2_RVT U1026 ( .A1(net31242), .A2(net31244), .A3(net48659), .Y(
        quotient[43]) );
  NAND4X0_RVT U1027 ( .A1(\u_div/CryTmp[43][4] ), .A2(net32156), .A3(net32118), 
        .A4(net31250), .Y(net31243) );
  INVX0_RVT U1028 ( .A(\u_div/SumTmp[43][2] ), .Y(n360) );
  INVX0_RVT U1029 ( .A(\u_div/SumTmp[43][1] ), .Y(n361) );
  INVX1_RVT U1030 ( .A(a[44]), .Y(n373) );
  XOR2X1_RVT U1031 ( .A1(a[44]), .A2(net32408), .Y(n374) );
  NOR3X2_RVT U1032 ( .A1(n363), .A2(n364), .A3(n376), .Y(quotient[44]) );
  NAND4X0_RVT U1033 ( .A1(n369), .A2(n370), .A3(n371), .A4(n372), .Y(n363) );
  NOR2X0_RVT U1034 ( .A1(net31872), .A2(net31896), .Y(n369) );
  INVX1_RVT U1035 ( .A(net31874), .Y(net31872) );
  INVX1_RVT U1036 ( .A(net31902), .Y(net31896) );
  NOR3X0_RVT U1037 ( .A1(net31844), .A2(net31814), .A3(net32352), .Y(n370) );
  INVX1_RVT U1038 ( .A(net31846), .Y(net31844) );
  INVX1_RVT U1039 ( .A(net31822), .Y(net31814) );
  INVX1_RVT U1040 ( .A(net32354), .Y(net32352) );
  NOR3X0_RVT U1041 ( .A1(net32300), .A2(net32264), .A3(net32324), .Y(n371) );
  INVX1_RVT U1042 ( .A(net32302), .Y(net32300) );
  INVX1_RVT U1043 ( .A(net32272), .Y(net32264) );
  INVX1_RVT U1044 ( .A(net32326), .Y(net32324) );
  NOR3X0_RVT U1045 ( .A1(net32234), .A2(net32210), .A3(net32178), .Y(n372) );
  INVX1_RVT U1046 ( .A(net32212), .Y(net32210) );
  INVX1_RVT U1047 ( .A(net32186), .Y(net32178) );
  NAND2X0_RVT U1048 ( .A1(n367), .A2(n368), .Y(n364) );
  NOR3X0_RVT U1049 ( .A1(net32024), .A2(b[14]), .A3(net31998), .Y(n367) );
  INVX1_RVT U1050 ( .A(net32032), .Y(net32024) );
  INVX1_RVT U1051 ( .A(net32002), .Y(net31998) );
  NOR3X0_RVT U1052 ( .A1(net31950), .A2(net31972), .A3(net31922), .Y(n368) );
  INVX1_RVT U1053 ( .A(net31952), .Y(net31950) );
  INVX1_RVT U1054 ( .A(net31930), .Y(net31922) );
  IBUFFX16_RVT U1055 ( .A(n365), .Y(n375) );
  NAND4X0_RVT U1056 ( .A1(\u_div/CryTmp[44][3] ), .A2(net32156), .A3(n366), 
        .A4(net32092), .Y(n365) );
  INVX1_RVT U1057 ( .A(n327), .Y(\u_div/PartRem[45][2] ) );
  MUX21X1_RVT U1058 ( .A1(net29755), .A2(net30099), .S0(quotient[45]), .Y(n327) );
  OR2X1_RVT U1059 ( .A1(net32408), .A2(a[44]), .Y(\u_div/CryTmp[44][1] ) );
  INVX2_RVT U1060 ( .A(n328), .Y(\u_div/PartRem[45][1] ) );
  MUX21X2_RVT U1061 ( .A1(net37220), .A2(net31434), .S0(net37219), .Y(n328) );
  INVX1_RVT U1062 ( .A(b[10]), .Y(net32156) );
  NOR2X0_RVT U1063 ( .A1(net32128), .A2(net32076), .Y(n366) );
  INVX1_RVT U1064 ( .A(net49055), .Y(net32128) );
  INVX1_RVT U1065 ( .A(net32078), .Y(net32076) );
  INVX1_RVT U1066 ( .A(net32104), .Y(net32092) );
  INVX0_RVT U1067 ( .A(\u_div/SumTmp[30][16] ), .Y(n424) );
  INVX1_RVT U1068 ( .A(n447), .Y(n448) );
  IBUFFX4_RVT U1069 ( .A(\u_div/CryTmp[30][16] ), .Y(n447) );
  MUX21X1_RVT U1070 ( .A1(net29900), .A2(net30148), .S0(net40084), .Y(n423) );
  INVX1_RVT U1071 ( .A(net32024), .Y(net32016) );
  MUX21X1_RVT U1072 ( .A1(net29901), .A2(net30208), .S0(net39869), .Y(net29916) );
  INVX1_RVT U1073 ( .A(b[14]), .Y(net32046) );
  INVX1_RVT U1074 ( .A(net29917), .Y(\u_div/PartRem[31][13] ) );
  MUX21X1_RVT U1075 ( .A1(net29902), .A2(net30256), .S0(net39874), .Y(net29917) );
  IBUFFX4_RVT U1076 ( .A(n449), .Y(n450) );
  IBUFFX4_RVT U1077 ( .A(\u_div/CryTmp[30][13] ), .Y(n442) );
  INVX1_RVT U1078 ( .A(net29918), .Y(\u_div/PartRem[31][12] ) );
  MUX21X1_RVT U1079 ( .A1(net29903), .A2(net30499), .S0(net39869), .Y(net29918) );
  INVX1_RVT U1080 ( .A(net32104), .Y(net32088) );
  INVX1_RVT U1081 ( .A(net29919), .Y(\u_div/PartRem[31][11] ) );
  MUX21X1_RVT U1082 ( .A1(net29904), .A2(net30547), .S0(net40084), .Y(net29919) );
  INVX1_RVT U1083 ( .A(net29920), .Y(\u_div/PartRem[31][10] ) );
  MUX21X1_RVT U1084 ( .A1(net29890), .A2(net30595), .S0(net39869), .Y(net29920) );
  INVX1_RVT U1085 ( .A(net32154), .Y(net32140) );
  INVX1_RVT U1086 ( .A(net29905), .Y(\u_div/PartRem[31][9] ) );
  MUX21X1_RVT U1087 ( .A1(net29891), .A2(net30643), .S0(net40084), .Y(net29905) );
  INVX1_RVT U1088 ( .A(net32178), .Y(net32166) );
  INVX1_RVT U1089 ( .A(net29906), .Y(\u_div/PartRem[31][8] ) );
  MUX21X1_RVT U1090 ( .A1(net29892), .A2(net30691), .S0(net39869), .Y(net29906) );
  INVX1_RVT U1091 ( .A(net32210), .Y(net32200) );
  INVX1_RVT U1092 ( .A(net29907), .Y(\u_div/PartRem[31][7] ) );
  MUX21X1_RVT U1093 ( .A1(net29893), .A2(net30739), .S0(net40084), .Y(net29907) );
  INVX1_RVT U1094 ( .A(net32234), .Y(net32222) );
  INVX1_RVT U1095 ( .A(net29908), .Y(\u_div/PartRem[31][6] ) );
  MUX21X1_RVT U1096 ( .A1(net29894), .A2(net30787), .S0(net39869), .Y(net29908) );
  INVX1_RVT U1097 ( .A(net32264), .Y(net32254) );
  IBUFFX16_RVT U1098 ( .A(net29909), .Y(\u_div/PartRem[31][5] ) );
  INVX1_RVT U1099 ( .A(net32300), .Y(net32284) );
  IBUFFX16_RVT U1100 ( .A(\u_div/CryTmp[30][5] ), .Y(n455) );
  INVX1_RVT U1101 ( .A(net29910), .Y(\u_div/PartRem[31][4] ) );
  MUX21X1_RVT U1102 ( .A1(net29896), .A2(net30883), .S0(net39869), .Y(net29910) );
  INVX1_RVT U1103 ( .A(net32324), .Y(net32314) );
  INVX1_RVT U1104 ( .A(net29911), .Y(\u_div/PartRem[31][3] ) );
  MUX21X1_RVT U1105 ( .A1(net29897), .A2(net30967), .S0(net40084), .Y(net29911) );
  INVX1_RVT U1106 ( .A(net32352), .Y(net32338) );
  IBUFFX16_RVT U1107 ( .A(\u_div/CryTmp[30][3] ), .Y(n453) );
  INVX1_RVT U1108 ( .A(net29912), .Y(\u_div/PartRem[31][2] ) );
  MUX21X2_RVT U1109 ( .A1(net29898), .A2(net30993), .S0(net40084), .Y(net29912) );
  INVX1_RVT U1110 ( .A(b[2]), .Y(net32366) );
  MUX21X1_RVT U1111 ( .A1(net31658), .A2(net37244), .S0(net39869), .Y(net29913) );
  INVX1_RVT U1112 ( .A(b[1]), .Y(net32386) );
  OR2X1_RVT U1113 ( .A1(net32406), .A2(a[30]), .Y(\u_div/CryTmp[30][1] ) );
  INVX1_RVT U1114 ( .A(net31998), .Y(net31982) );
  IBUFFX32_RVT U1115 ( .A(n422), .Y(\u_div/PartRem[31][16] ) );
  MUX21X1_RVT U1116 ( .A1(net29899), .A2(net30085), .S0(net40084), .Y(n422) );
  MUX21X1_RVT U1117 ( .A1(n422), .A2(n424), .S0(net37577), .Y(net29930) );
  IBUFFX16_RVT U1118 ( .A(\u_div/CryTmp[30][17] ), .Y(net31303) );
  INVX0_RVT U1119 ( .A(\u_div/SumTmp[30][15] ), .Y(net30147) );
  INVX1_RVT U1120 ( .A(net29900), .Y(\u_div/PartRem[32][14] ) );
  INVX1_RVT U1121 ( .A(net29901), .Y(\u_div/PartRem[32][13] ) );
  INVX1_RVT U1122 ( .A(net29902), .Y(\u_div/PartRem[32][12] ) );
  MUX21X1_RVT U1123 ( .A1(n420), .A2(n427), .S0(net50050), .Y(net29902) );
  INVX1_RVT U1124 ( .A(net29903), .Y(\u_div/PartRem[32][11] ) );
  MUX21X1_RVT U1125 ( .A1(n421), .A2(net30500), .S0(net50049), .Y(net29903) );
  INVX1_RVT U1126 ( .A(net29904), .Y(\u_div/PartRem[32][10] ) );
  MUX21X1_RVT U1127 ( .A1(n409), .A2(net30548), .S0(net50050), .Y(net29904) );
  INVX1_RVT U1128 ( .A(net29890), .Y(\u_div/PartRem[32][9] ) );
  MUX21X1_RVT U1129 ( .A1(n410), .A2(net30596), .S0(net50049), .Y(net29890) );
  INVX1_RVT U1130 ( .A(net29891), .Y(\u_div/PartRem[32][8] ) );
  MUX21X1_RVT U1131 ( .A1(n411), .A2(net30644), .S0(net50050), .Y(net29891) );
  INVX4_RVT U1132 ( .A(n436), .Y(n437) );
  INVX1_RVT U1133 ( .A(net29892), .Y(\u_div/PartRem[32][7] ) );
  MUX21X1_RVT U1134 ( .A1(n412), .A2(net30692), .S0(net50049), .Y(net29892) );
  INVX1_RVT U1135 ( .A(net32234), .Y(net32226) );
  INVX1_RVT U1136 ( .A(net29893), .Y(\u_div/PartRem[32][6] ) );
  MUX21X1_RVT U1137 ( .A1(n413), .A2(net30740), .S0(net50050), .Y(net29893) );
  INVX1_RVT U1138 ( .A(net29894), .Y(\u_div/PartRem[32][5] ) );
  MUX21X1_RVT U1139 ( .A1(n414), .A2(net30788), .S0(net50049), .Y(net29894) );
  INVX1_RVT U1140 ( .A(net29895), .Y(\u_div/PartRem[32][4] ) );
  MUX21X1_RVT U1141 ( .A1(n415), .A2(net30836), .S0(net50050), .Y(net29895) );
  INVX1_RVT U1142 ( .A(net29896), .Y(\u_div/PartRem[32][3] ) );
  INVX1_RVT U1143 ( .A(net29897), .Y(\u_div/PartRem[32][2] ) );
  OR2X1_RVT U1144 ( .A1(net32406), .A2(a[31]), .Y(\u_div/CryTmp[31][1] ) );
  NBUFFX2_RVT U1145 ( .A(net39874), .Y(net40084) );
  MUX21X1_RVT U1146 ( .A1(n423), .A2(net30147), .S0(net37577), .Y(net29931) );
  MUX21X1_RVT U1147 ( .A1(net29873), .A2(net30150), .S0(net37854), .Y(n418) );
  INVX0_RVT U1148 ( .A(\u_div/SumTmp[32][13] ), .Y(n425) );
  IBUFFX4_RVT U1149 ( .A(n419), .Y(\u_div/PartRem[33][12] ) );
  MUX21X1_RVT U1150 ( .A1(net29874), .A2(net30210), .S0(net37854), .Y(n419) );
  INVX1_RVT U1151 ( .A(n420), .Y(\u_div/PartRem[33][11] ) );
  MUX21X1_RVT U1152 ( .A1(n408), .A2(n428), .S0(net37854), .Y(n420) );
  IBUFFX4_RVT U1153 ( .A(\u_div/CryTmp[32][11] ), .Y(n444) );
  INVX1_RVT U1154 ( .A(n421), .Y(\u_div/PartRem[33][10] ) );
  MUX21X1_RVT U1155 ( .A1(n399), .A2(n29), .S0(net37854), .Y(n421) );
  INVX1_RVT U1156 ( .A(n409), .Y(\u_div/PartRem[33][9] ) );
  MUX21X1_RVT U1157 ( .A1(n400), .A2(net30549), .S0(net37854), .Y(n409) );
  INVX1_RVT U1158 ( .A(n410), .Y(\u_div/PartRem[33][8] ) );
  MUX21X1_RVT U1159 ( .A1(net46421), .A2(net30597), .S0(net37854), .Y(n410) );
  INVX1_RVT U1160 ( .A(n411), .Y(\u_div/PartRem[33][7] ) );
  MUX21X1_RVT U1161 ( .A1(n402), .A2(net30645), .S0(net37854), .Y(n411) );
  INVX1_RVT U1162 ( .A(n412), .Y(\u_div/PartRem[33][6] ) );
  MUX21X1_RVT U1163 ( .A1(n403), .A2(net30693), .S0(net37854), .Y(n412) );
  INVX1_RVT U1164 ( .A(n413), .Y(\u_div/PartRem[33][5] ) );
  MUX21X1_RVT U1165 ( .A1(n404), .A2(net30741), .S0(net37854), .Y(n413) );
  INVX1_RVT U1166 ( .A(n414), .Y(\u_div/PartRem[33][4] ) );
  MUX21X1_RVT U1167 ( .A1(n405), .A2(net30789), .S0(net37854), .Y(n414) );
  INVX1_RVT U1168 ( .A(n415), .Y(\u_div/PartRem[33][3] ) );
  MUX21X1_RVT U1169 ( .A1(n406), .A2(net30837), .S0(net37854), .Y(n415) );
  INVX1_RVT U1170 ( .A(n416), .Y(\u_div/PartRem[33][2] ) );
  MUX21X1_RVT U1171 ( .A1(n407), .A2(net30885), .S0(net37854), .Y(n416) );
  INVX1_RVT U1172 ( .A(n417), .Y(\u_div/PartRem[33][1] ) );
  MUX21X1_RVT U1173 ( .A1(net31626), .A2(net37231), .S0(net37854), .Y(n417) );
  OR2X1_RVT U1174 ( .A1(net32406), .A2(a[32]), .Y(\u_div/CryTmp[32][1] ) );
  NOR2X2_RVT U1175 ( .A1(net31297), .A2(n434), .Y(net50049) );
  OR2X1_RVT U1176 ( .A1(net31998), .A2(net31295), .Y(net31297) );
  NAND2X0_RVT U1177 ( .A1(net52311), .A2(\u_div/CryTmp[32][15] ), .Y(n434) );
  INVX1_RVT U1178 ( .A(net29885), .Y(\u_div/PartRem[33][14] ) );
  MUX21X1_RVT U1179 ( .A1(net29872), .A2(net30087), .S0(net37854), .Y(net29885) );
  NOR2X1_RVT U1180 ( .A1(net31297), .A2(n434), .Y(n435) );
  NOR2X2_RVT U1181 ( .A1(net31297), .A2(n434), .Y(net50050) );
  INVX0_RVT U1182 ( .A(\u_div/SumTmp[32][14] ), .Y(net30086) );
  INVX0_RVT U1183 ( .A(\u_div/SumTmp[32][11] ), .Y(n427) );
  IBUFFX16_RVT U1184 ( .A(\u_div/SumTmp[33][10] ), .Y(n428) );
  INVX0_RVT U1185 ( .A(n408), .Y(\u_div/PartRem[34][10] ) );
  INVX1_RVT U1186 ( .A(n399), .Y(\u_div/PartRem[34][9] ) );
  MUX21X1_RVT U1187 ( .A1(net46238), .A2(n429), .S0(net37563), .Y(n399) );
  INVX1_RVT U1188 ( .A(n400), .Y(\u_div/PartRem[34][8] ) );
  MUX21X1_RVT U1189 ( .A1(n393), .A2(n430), .S0(net37563), .Y(n400) );
  MUX21X1_RVT U1190 ( .A1(net29854), .A2(net30598), .S0(net37563), .Y(n401) );
  MUX21X1_RVT U1191 ( .A1(net29844), .A2(net30599), .S0(net50471), .Y(net29854) );
  IBUFFX16_RVT U1192 ( .A(\u_div/SumTmp[34][6] ), .Y(net30598) );
  INVX1_RVT U1193 ( .A(n402), .Y(\u_div/PartRem[34][6] ) );
  MUX21X1_RVT U1194 ( .A1(n394), .A2(n431), .S0(net37563), .Y(n402) );
  INVX1_RVT U1195 ( .A(n403), .Y(\u_div/PartRem[34][5] ) );
  MUX21X1_RVT U1196 ( .A1(n395), .A2(net30694), .S0(net37563), .Y(n403) );
  INVX1_RVT U1197 ( .A(n404), .Y(\u_div/PartRem[34][4] ) );
  MUX21X1_RVT U1198 ( .A1(n396), .A2(net30742), .S0(net37563), .Y(n404) );
  INVX1_RVT U1199 ( .A(n405), .Y(\u_div/PartRem[34][3] ) );
  MUX21X1_RVT U1200 ( .A1(n397), .A2(net30790), .S0(net37563), .Y(n405) );
  INVX1_RVT U1201 ( .A(n406), .Y(\u_div/PartRem[34][2] ) );
  MUX21X1_RVT U1202 ( .A1(n398), .A2(net30838), .S0(net37563), .Y(n406) );
  INVX1_RVT U1203 ( .A(n407), .Y(\u_div/PartRem[34][1] ) );
  MUX21X1_RVT U1204 ( .A1(net31610), .A2(net37246), .S0(net37563), .Y(n407) );
  OR2X1_RVT U1205 ( .A1(net32406), .A2(a[33]), .Y(\u_div/CryTmp[33][1] ) );
  NOR2X4_RVT U1206 ( .A1(net31292), .A2(net31294), .Y(net37854) );
  INVX16_RVT U1207 ( .A(n278), .Y(\u_div/PartRem[35][9] ) );
  INVX1_RVT U1208 ( .A(n393), .Y(\u_div/PartRem[35][7] ) );
  MUX21X1_RVT U1209 ( .A1(net29843), .A2(net30551), .S0(net50471), .Y(n393) );
  INVX1_RVT U1210 ( .A(net29854), .Y(\u_div/PartRem[35][6] ) );
  MUX21X1_RVT U1211 ( .A1(n389), .A2(n432), .S0(net50471), .Y(n394) );
  INVX1_RVT U1212 ( .A(n395), .Y(\u_div/PartRem[35][4] ) );
  MUX21X1_RVT U1213 ( .A1(net52890), .A2(net30695), .S0(net50471), .Y(n395) );
  INVX1_RVT U1214 ( .A(n396), .Y(\u_div/PartRem[35][3] ) );
  MUX21X1_RVT U1215 ( .A1(n390), .A2(net30743), .S0(net50471), .Y(n396) );
  INVX1_RVT U1216 ( .A(n397), .Y(\u_div/PartRem[35][2] ) );
  MUX21X1_RVT U1217 ( .A1(n391), .A2(net30791), .S0(net50471), .Y(n397) );
  MUX21X1_RVT U1218 ( .A1(net31594), .A2(net37247), .S0(net50471), .Y(n398) );
  OR2X1_RVT U1219 ( .A1(net32406), .A2(a[34]), .Y(\u_div/CryTmp[34][1] ) );
  INVX0_RVT U1220 ( .A(\u_div/SumTmp[34][7] ), .Y(n430) );
  IBUFFX16_RVT U1221 ( .A(\u_div/SumTmp[34][5] ), .Y(n431) );
  MUX21X1_RVT U1222 ( .A1(net29836), .A2(n433), .S0(net37570), .Y(n389) );
  INVX0_RVT U1223 ( .A(\u_div/SumTmp[35][4] ), .Y(n432) );
  IBUFFX4_RVT U1224 ( .A(n389), .Y(\u_div/PartRem[36][4] ) );
  IBUFFX4_RVT U1225 ( .A(net29846), .Y(\u_div/PartRem[36][3] ) );
  INVX1_RVT U1226 ( .A(n390), .Y(\u_div/PartRem[36][2] ) );
  MUX21X1_RVT U1227 ( .A1(n388), .A2(net30744), .S0(net37570), .Y(n390) );
  INVX1_RVT U1228 ( .A(n391), .Y(\u_div/PartRem[36][1] ) );
  MUX21X1_RVT U1229 ( .A1(net31578), .A2(net37251), .S0(net37570), .Y(n391) );
  OR2X1_RVT U1230 ( .A1(net32406), .A2(a[35]), .Y(\u_div/CryTmp[35][1] ) );
  INVX4_RVT U1231 ( .A(net50470), .Y(net50471) );
  INVX0_RVT U1232 ( .A(\u_div/SumTmp[36][3] ), .Y(n433) );
  IBUFFX16_RVT U1233 ( .A(net29836), .Y(\u_div/PartRem[37][3] ) );
  IBUFFX16_RVT U1234 ( .A(net29837), .Y(\u_div/PartRem[37][2] ) );
  IBUFFX16_RVT U1235 ( .A(n388), .Y(\u_div/PartRem[37][1] ) );
  MUX21X2_RVT U1236 ( .A1(net31562), .A2(net37249), .S0(net37242), .Y(n388) );
  OR2X1_RVT U1237 ( .A1(net32408), .A2(a[36]), .Y(\u_div/CryTmp[36][1] ) );
  NOR2X2_RVT U1238 ( .A1(net31255), .A2(net31281), .Y(net37570) );
  INVX1_RVT U1239 ( .A(net46015), .Y(net29828) );
  NOR2X2_RVT U1240 ( .A1(b[10]), .A2(net43355), .Y(net37242) );
  MUX21X1_RVT U1241 ( .A1(net29974), .A2(net30081), .S0(net41415), .Y(net29992) );
  INVX1_RVT U1242 ( .A(net31896), .Y(net31882) );
  INVX1_RVT U1243 ( .A(net29994), .Y(\u_div/PartRem[27][19] ) );
  INVX1_RVT U1244 ( .A(net31922), .Y(net31914) );
  INVX1_RVT U1245 ( .A(net29995), .Y(\u_div/PartRem[27][18] ) );
  MUX21X1_RVT U1246 ( .A1(net29976), .A2(net30204), .S0(net41415), .Y(net29995) );
  INVX1_RVT U1247 ( .A(net31950), .Y(net31938) );
  INVX1_RVT U1248 ( .A(net29996), .Y(\u_div/PartRem[27][17] ) );
  MUX21X1_RVT U1249 ( .A1(net29977), .A2(net30252), .S0(net41415), .Y(net29996) );
  INVX1_RVT U1250 ( .A(net31972), .Y(net31960) );
  INVX1_RVT U1251 ( .A(net29997), .Y(\u_div/PartRem[27][16] ) );
  MUX21X1_RVT U1252 ( .A1(net29978), .A2(net30495), .S0(net41415), .Y(net29997) );
  INVX0_RVT U1253 ( .A(net29998), .Y(\u_div/PartRem[27][15] ) );
  MUX21X1_RVT U1254 ( .A1(net29979), .A2(net30543), .S0(net41415), .Y(net29998) );
  INVX1_RVT U1255 ( .A(net29999), .Y(\u_div/PartRem[27][14] ) );
  MUX21X1_RVT U1256 ( .A1(net29980), .A2(net30591), .S0(net41415), .Y(net29999) );
  MUX21X1_RVT U1257 ( .A1(net29981), .A2(net30639), .S0(net41415), .Y(net30000) );
  INVX1_RVT U1258 ( .A(net30001), .Y(\u_div/PartRem[27][12] ) );
  MUX21X1_RVT U1259 ( .A1(net29982), .A2(net49675), .S0(net41415), .Y(net30001) );
  MUX21X1_RVT U1260 ( .A1(net29965), .A2(net30783), .S0(net41415), .Y(net30003) );
  INVX1_RVT U1261 ( .A(net29984), .Y(\u_div/PartRem[27][9] ) );
  MUX21X1_RVT U1262 ( .A1(net29966), .A2(net30831), .S0(net41415), .Y(net29984) );
  INVX1_RVT U1263 ( .A(net32178), .Y(net32168) );
  INVX1_RVT U1264 ( .A(net29985), .Y(\u_div/PartRem[27][8] ) );
  MUX21X1_RVT U1265 ( .A1(net29967), .A2(net30879), .S0(net41415), .Y(net29985) );
  INVX1_RVT U1266 ( .A(net29986), .Y(\u_div/PartRem[27][7] ) );
  INVX1_RVT U1267 ( .A(net29987), .Y(\u_div/PartRem[27][6] ) );
  MUX21X1_RVT U1268 ( .A1(net29969), .A2(net30989), .S0(net41415), .Y(net29987) );
  INVX1_RVT U1269 ( .A(net29989), .Y(\u_div/PartRem[27][4] ) );
  MUX21X1_RVT U1270 ( .A1(net29971), .A2(net31036), .S0(net41415), .Y(net29989) );
  INVX1_RVT U1271 ( .A(net29990), .Y(\u_div/PartRem[27][3] ) );
  MUX21X1_RVT U1272 ( .A1(net29972), .A2(net31058), .S0(net41415), .Y(net29990) );
  INVX1_RVT U1273 ( .A(net29991), .Y(\u_div/PartRem[27][2] ) );
  MUX21X1_RVT U1274 ( .A1(net29973), .A2(net31080), .S0(net41415), .Y(net29991) );
  INVX1_RVT U1275 ( .A(net29993), .Y(\u_div/PartRem[27][1] ) );
  MUX21X1_RVT U1276 ( .A1(net31722), .A2(net37248), .S0(net41415), .Y(net29993) );
  OR2X1_RVT U1277 ( .A1(net32406), .A2(a[26]), .Y(\u_div/CryTmp[26][1] ) );
  INVX1_RVT U1278 ( .A(net29988), .Y(\u_div/PartRem[27][5] ) );
  MUX21X1_RVT U1279 ( .A1(net29970), .A2(net31013), .S0(net41415), .Y(net29988) );
  MUX21X1_RVT U1280 ( .A1(net29983), .A2(net49672), .S0(net41415), .Y(net30002) );
  INVX0_RVT U1281 ( .A(\u_div/SumTmp[26][20] ), .Y(net30080) );
  INVX0_RVT U1282 ( .A(\u_div/SumTmp[26][19] ), .Y(net30143) );
  IBUFFX16_RVT U1283 ( .A(\u_div/SumTmp[26][18] ), .Y(net30203) );
  INVX0_RVT U1284 ( .A(\u_div/SumTmp[26][17] ), .Y(net30251) );
  INVX0_RVT U1285 ( .A(\u_div/SumTmp[26][16] ), .Y(net30494) );
  INVX0_RVT U1286 ( .A(\u_div/SumTmp[26][15] ), .Y(net30542) );
  INVX0_RVT U1287 ( .A(\u_div/SumTmp[26][14] ), .Y(net30590) );
  INVX0_RVT U1288 ( .A(\u_div/SumTmp[26][13] ), .Y(net30638) );
  INVX0_RVT U1289 ( .A(\u_div/SumTmp[26][12] ), .Y(net30686) );
  INVX0_RVT U1290 ( .A(\u_div/SumTmp[26][11] ), .Y(net30734) );
  MUX21X1_RVT U1291 ( .A1(n465), .A2(n475), .S0(quotient[28]), .Y(net29983) );
  NBUFFX8_RVT U1292 ( .A(net30735), .Y(net49672) );
  INVX1_RVT U1293 ( .A(net32154), .Y(net32142) );
  INVX1_RVT U1294 ( .A(net29965), .Y(\u_div/PartRem[28][9] ) );
  MUX21X1_RVT U1295 ( .A1(n466), .A2(n476), .S0(quotient[28]), .Y(net29965) );
  MUX21X1_RVT U1296 ( .A1(n467), .A2(n477), .S0(quotient[28]), .Y(net29966) );
  INVX1_RVT U1297 ( .A(net29967), .Y(\u_div/PartRem[28][7] ) );
  MUX21X1_RVT U1298 ( .A1(n468), .A2(n478), .S0(quotient[28]), .Y(net29967) );
  INVX1_RVT U1299 ( .A(net29968), .Y(\u_div/PartRem[28][6] ) );
  MUX21X1_RVT U1300 ( .A1(n469), .A2(n479), .S0(quotient[28]), .Y(net29968) );
  INVX1_RVT U1301 ( .A(net29969), .Y(\u_div/PartRem[28][5] ) );
  MUX21X1_RVT U1302 ( .A1(n470), .A2(n480), .S0(quotient[28]), .Y(net29969) );
  INVX1_RVT U1303 ( .A(net29970), .Y(\u_div/PartRem[28][4] ) );
  MUX21X1_RVT U1304 ( .A1(n471), .A2(n481), .S0(quotient[28]), .Y(net29970) );
  MUX21X1_RVT U1305 ( .A1(n472), .A2(n482), .S0(quotient[28]), .Y(net29971) );
  IBUFFX16_RVT U1306 ( .A(\u_div/CryTmp[27][3] ), .Y(n487) );
  INVX1_RVT U1307 ( .A(net29972), .Y(\u_div/PartRem[28][2] ) );
  MUX21X1_RVT U1308 ( .A1(n473), .A2(n483), .S0(quotient[28]), .Y(net29972) );
  INVX1_RVT U1309 ( .A(net29973), .Y(\u_div/PartRem[28][1] ) );
  MUX21X1_RVT U1310 ( .A1(net31706), .A2(net37263), .S0(quotient[28]), .Y(
        net29973) );
  OR2X1_RVT U1311 ( .A1(net32406), .A2(a[27]), .Y(\u_div/CryTmp[27][1] ) );
  AND2X1_RVT U1312 ( .A1(net31272), .A2(\u_div/CryTmp[27][20] ), .Y(net41415)
         );
  MUX21X1_RVT U1313 ( .A1(n457), .A2(net30737), .S0(net47679), .Y(n465) );
  INVX0_RVT U1314 ( .A(\u_div/SumTmp[28][9] ), .Y(n475) );
  INVX1_RVT U1315 ( .A(n465), .Y(\u_div/PartRem[29][9] ) );
  INVX1_RVT U1316 ( .A(n466), .Y(\u_div/PartRem[29][8] ) );
  MUX21X1_RVT U1317 ( .A1(n458), .A2(net30785), .S0(net47679), .Y(n466) );
  INVX1_RVT U1318 ( .A(n467), .Y(\u_div/PartRem[29][7] ) );
  MUX21X1_RVT U1319 ( .A1(n459), .A2(net30833), .S0(net47679), .Y(n467) );
  INVX1_RVT U1320 ( .A(net32234), .Y(net32224) );
  INVX1_RVT U1321 ( .A(n468), .Y(\u_div/PartRem[29][6] ) );
  MUX21X1_RVT U1322 ( .A1(n460), .A2(net30881), .S0(net47679), .Y(n468) );
  INVX1_RVT U1323 ( .A(n469), .Y(\u_div/PartRem[29][5] ) );
  MUX21X1_RVT U1324 ( .A1(n461), .A2(net30965), .S0(net47679), .Y(n469) );
  INVX1_RVT U1325 ( .A(n470), .Y(\u_div/PartRem[29][4] ) );
  MUX21X1_RVT U1326 ( .A1(n462), .A2(net30991), .S0(net47679), .Y(n470) );
  INVX1_RVT U1327 ( .A(n471), .Y(\u_div/PartRem[29][3] ) );
  MUX21X1_RVT U1328 ( .A1(n463), .A2(net31015), .S0(net47679), .Y(n471) );
  INVX1_RVT U1329 ( .A(n472), .Y(\u_div/PartRem[29][2] ) );
  MUX21X1_RVT U1330 ( .A1(n464), .A2(net31038), .S0(net47679), .Y(n472) );
  OR2X1_RVT U1331 ( .A1(net32406), .A2(a[28]), .Y(\u_div/CryTmp[28][1] ) );
  INVX1_RVT U1332 ( .A(n473), .Y(\u_div/PartRem[29][1] ) );
  MUX21X1_RVT U1333 ( .A1(n485), .A2(n486), .S0(net47679), .Y(n473) );
  INVX2_RVT U1334 ( .A(net31310), .Y(quotient[28]) );
  IBUFFX16_RVT U1335 ( .A(\u_div/CryTmp[28][10] ), .Y(net42938) );
  IBUFFX16_RVT U1336 ( .A(\u_div/SumTmp[28][8] ), .Y(n476) );
  IBUFFX16_RVT U1337 ( .A(\u_div/SumTmp[28][7] ), .Y(n477) );
  INVX0_RVT U1338 ( .A(\u_div/SumTmp[28][6] ), .Y(n478) );
  INVX0_RVT U1339 ( .A(\u_div/SumTmp[28][5] ), .Y(n479) );
  INVX0_RVT U1340 ( .A(\u_div/SumTmp[28][4] ), .Y(n480) );
  INVX0_RVT U1341 ( .A(\u_div/SumTmp[28][3] ), .Y(n481) );
  INVX0_RVT U1342 ( .A(\u_div/SumTmp[28][2] ), .Y(n482) );
  INVX0_RVT U1343 ( .A(\u_div/SumTmp[28][1] ), .Y(n483) );
  INVX1_RVT U1344 ( .A(a[29]), .Y(n485) );
  XOR2X1_RVT U1345 ( .A1(a[29]), .A2(net32406), .Y(n486) );
  NOR2X1_RVT U1346 ( .A1(net31922), .A2(net31276), .Y(net47690) );
  INVX1_RVT U1347 ( .A(net29930), .Y(\u_div/PartRem[30][17] ) );
  INVX1_RVT U1348 ( .A(net29931), .Y(\u_div/PartRem[30][16] ) );
  INVX4_RVT U1349 ( .A(n497), .Y(n498) );
  INVX4_RVT U1350 ( .A(n490), .Y(n497) );
  IBUFFX16_RVT U1351 ( .A(n489), .Y(n490) );
  INVX32_RVT U1352 ( .A(\u_div/CryTmp[29][16] ), .Y(n489) );
  INVX1_RVT U1353 ( .A(net29932), .Y(\u_div/PartRem[30][15] ) );
  MUX21X1_RVT U1354 ( .A1(net29916), .A2(net30207), .S0(net37577), .Y(net29932) );
  INVX1_RVT U1355 ( .A(net29933), .Y(\u_div/PartRem[30][14] ) );
  MUX21X1_RVT U1356 ( .A1(net29917), .A2(net30255), .S0(net37577), .Y(net29933) );
  MUX21X1_RVT U1357 ( .A1(net29918), .A2(net30498), .S0(net37577), .Y(net29934) );
  INVX1_RVT U1358 ( .A(net29935), .Y(\u_div/PartRem[30][12] ) );
  MUX21X1_RVT U1359 ( .A1(net29919), .A2(net30546), .S0(net37577), .Y(net29935) );
  INVX1_RVT U1360 ( .A(net29936), .Y(\u_div/PartRem[30][11] ) );
  MUX21X1_RVT U1361 ( .A1(net29920), .A2(net30594), .S0(net37577), .Y(net29936) );
  INVX1_RVT U1362 ( .A(net29937), .Y(\u_div/PartRem[30][10] ) );
  MUX21X1_RVT U1363 ( .A1(net29905), .A2(net30642), .S0(net37577), .Y(net29937) );
  INVX1_RVT U1364 ( .A(net29921), .Y(\u_div/PartRem[30][9] ) );
  MUX21X1_RVT U1365 ( .A1(net29906), .A2(net30690), .S0(net37577), .Y(net29921) );
  INVX1_RVT U1366 ( .A(n458), .Y(\u_div/PartRem[30][7] ) );
  MUX21X1_RVT U1367 ( .A1(net29908), .A2(net30786), .S0(net37577), .Y(n458) );
  INVX1_RVT U1368 ( .A(n459), .Y(\u_div/PartRem[30][6] ) );
  MUX21X1_RVT U1369 ( .A1(net29909), .A2(net30834), .S0(net37577), .Y(n459) );
  INVX1_RVT U1370 ( .A(n460), .Y(\u_div/PartRem[30][5] ) );
  MUX21X1_RVT U1371 ( .A1(net29910), .A2(net30882), .S0(net37577), .Y(n460) );
  INVX1_RVT U1372 ( .A(n461), .Y(\u_div/PartRem[30][4] ) );
  MUX21X1_RVT U1373 ( .A1(net29911), .A2(net30966), .S0(net37577), .Y(n461) );
  INVX1_RVT U1374 ( .A(n462), .Y(\u_div/PartRem[30][3] ) );
  MUX21X1_RVT U1375 ( .A1(net29912), .A2(net52536), .S0(net37577), .Y(n462) );
  INVX1_RVT U1376 ( .A(n463), .Y(\u_div/PartRem[30][2] ) );
  MUX21X1_RVT U1377 ( .A1(net29913), .A2(net52534), .S0(net37577), .Y(n463) );
  INVX1_RVT U1378 ( .A(n464), .Y(\u_div/PartRem[30][1] ) );
  OR2X1_RVT U1379 ( .A1(net32406), .A2(a[29]), .Y(\u_div/CryTmp[29][1] ) );
  INVX0_RVT U1380 ( .A(\u_div/SumTmp[29][17] ), .Y(n474) );
  NOR2X4_RVT U1381 ( .A1(net31295), .A2(net52520), .Y(net37577) );
  MUX21X1_RVT U1382 ( .A1(net29930), .A2(n474), .S0(net47679), .Y(net29956) );
  INVX1_RVT U1383 ( .A(net30037), .Y(\u_div/PartRem[25][19] ) );
  MUX21X1_RVT U1384 ( .A1(net30016), .A2(net30250), .S0(quotient[25]), .Y(
        net30037) );
  INVX1_RVT U1385 ( .A(net30038), .Y(\u_div/PartRem[25][18] ) );
  MUX21X1_RVT U1386 ( .A1(net30017), .A2(net30493), .S0(quotient[25]), .Y(
        net30038) );
  INVX1_RVT U1387 ( .A(net30039), .Y(\u_div/PartRem[25][17] ) );
  MUX21X1_RVT U1388 ( .A1(net30018), .A2(net30541), .S0(quotient[25]), .Y(
        net30039) );
  INVX1_RVT U1389 ( .A(net30040), .Y(\u_div/PartRem[25][16] ) );
  MUX21X1_RVT U1390 ( .A1(net30019), .A2(net30589), .S0(quotient[25]), .Y(
        net30040) );
  INVX1_RVT U1391 ( .A(net30041), .Y(\u_div/PartRem[25][15] ) );
  MUX21X1_RVT U1392 ( .A1(net30020), .A2(net30637), .S0(quotient[25]), .Y(
        net30041) );
  INVX1_RVT U1393 ( .A(n499), .Y(\u_div/PartRem[25][14] ) );
  INVX1_RVT U1394 ( .A(n500), .Y(\u_div/PartRem[25][13] ) );
  MUX21X1_RVT U1395 ( .A1(net30022), .A2(net30733), .S0(quotient[25]), .Y(n500) );
  INVX1_RVT U1396 ( .A(\u_div/SumTmp[25][12] ), .Y(net30733) );
  INVX8_RVT U1397 ( .A(net31317), .Y(quotient[25]) );
  IBUFFX16_RVT U1398 ( .A(\u_div/CryTmp[24][13] ), .Y(n513) );
  INVX1_RVT U1399 ( .A(net30044), .Y(\u_div/PartRem[25][12] ) );
  MUX21X1_RVT U1400 ( .A1(net30023), .A2(net30781), .S0(quotient[25]), .Y(
        net30044) );
  INVX1_RVT U1401 ( .A(net30045), .Y(\u_div/PartRem[25][11] ) );
  MUX21X1_RVT U1402 ( .A1(net30024), .A2(net30829), .S0(quotient[25]), .Y(
        net30045) );
  INVX1_RVT U1403 ( .A(n501), .Y(\u_div/PartRem[25][10] ) );
  MUX21X1_RVT U1404 ( .A1(net29985), .A2(net30878), .S0(n145), .Y(net30004) );
  IBUFFX16_RVT U1405 ( .A(\u_div/SumTmp[25][9] ), .Y(net30877) );
  INVX1_RVT U1406 ( .A(net30025), .Y(\u_div/PartRem[25][9] ) );
  MUX21X1_RVT U1407 ( .A1(net30005), .A2(net30961), .S0(quotient[25]), .Y(
        net30025) );
  INVX1_RVT U1408 ( .A(net30026), .Y(\u_div/PartRem[25][8] ) );
  MUX21X1_RVT U1409 ( .A1(net30006), .A2(net30987), .S0(quotient[25]), .Y(
        net30026) );
  INVX1_RVT U1410 ( .A(net30027), .Y(\u_div/PartRem[25][7] ) );
  MUX21X1_RVT U1411 ( .A1(net30007), .A2(net31011), .S0(quotient[25]), .Y(
        net30027) );
  INVX1_RVT U1412 ( .A(net30028), .Y(\u_div/PartRem[25][6] ) );
  MUX21X1_RVT U1413 ( .A1(net30008), .A2(net31034), .S0(quotient[25]), .Y(
        net30028) );
  INVX1_RVT U1414 ( .A(net30029), .Y(\u_div/PartRem[25][5] ) );
  MUX21X1_RVT U1415 ( .A1(net30009), .A2(n91), .S0(quotient[25]), .Y(net30029)
         );
  INVX4_RVT U1416 ( .A(n507), .Y(n508) );
  IBUFFX16_RVT U1417 ( .A(\u_div/CryTmp[24][5] ), .Y(n507) );
  INVX1_RVT U1418 ( .A(net30030), .Y(\u_div/PartRem[25][4] ) );
  MUX21X1_RVT U1419 ( .A1(net30010), .A2(net31078), .S0(quotient[25]), .Y(
        net30030) );
  INVX1_RVT U1420 ( .A(net30031), .Y(\u_div/PartRem[25][3] ) );
  MUX21X1_RVT U1421 ( .A1(net30011), .A2(net31098), .S0(quotient[25]), .Y(
        net30031) );
  INVX1_RVT U1422 ( .A(net30032), .Y(\u_div/PartRem[25][2] ) );
  MUX21X1_RVT U1423 ( .A1(net30014), .A2(net31117), .S0(quotient[25]), .Y(
        net30032) );
  MUX21X2_RVT U1424 ( .A1(net41046), .A2(a[25]), .S0(net31317), .Y(net41045)
         );
  OR2X1_RVT U1425 ( .A1(net32406), .A2(a[24]), .Y(\u_div/CryTmp[24][1] ) );
  INVX0_RVT U1426 ( .A(\u_div/SumTmp[24][19] ), .Y(net30249) );
  INVX0_RVT U1427 ( .A(\u_div/SumTmp[24][18] ), .Y(net30492) );
  INVX0_RVT U1428 ( .A(\u_div/SumTmp[24][17] ), .Y(net30540) );
  INVX0_RVT U1429 ( .A(\u_div/SumTmp[24][16] ), .Y(net30588) );
  INVX0_RVT U1430 ( .A(\u_div/SumTmp[24][15] ), .Y(net30636) );
  INVX0_RVT U1431 ( .A(\u_div/SumTmp[24][14] ), .Y(net30684) );
  MUX21X1_RVT U1432 ( .A1(net30001), .A2(net30686), .S0(quotient[26]), .Y(
        net30021) );
  IBUFFX16_RVT U1433 ( .A(\u_div/SumTmp[25][13] ), .Y(net30685) );
  INVX1_RVT U1434 ( .A(net30022), .Y(\u_div/PartRem[26][12] ) );
  INVX1_RVT U1435 ( .A(net30023), .Y(\u_div/PartRem[26][11] ) );
  MUX21X1_RVT U1436 ( .A1(net30003), .A2(net30782), .S0(n153), .Y(net30023) );
  INVX1_RVT U1437 ( .A(net30024), .Y(\u_div/PartRem[26][10] ) );
  MUX21X1_RVT U1438 ( .A1(net29984), .A2(net30830), .S0(n144), .Y(net30024) );
  INVX1_RVT U1439 ( .A(net30004), .Y(\u_div/PartRem[26][9] ) );
  MUX21X1_RVT U1440 ( .A1(net29987), .A2(net30988), .S0(n145), .Y(net30006) );
  IBUFFX16_RVT U1441 ( .A(\u_div/CryTmp[25][7] ), .Y(n511) );
  INVX1_RVT U1442 ( .A(net30007), .Y(\u_div/PartRem[26][6] ) );
  MUX21X1_RVT U1443 ( .A1(net29988), .A2(net31012), .S0(n151), .Y(net30007) );
  INVX1_RVT U1444 ( .A(net30008), .Y(\u_div/PartRem[26][5] ) );
  MUX21X1_RVT U1445 ( .A1(net29989), .A2(net31035), .S0(n149), .Y(net30008) );
  INVX1_RVT U1446 ( .A(net30009), .Y(\u_div/PartRem[26][4] ) );
  MUX21X1_RVT U1447 ( .A1(net29990), .A2(net31057), .S0(n148), .Y(net30009) );
  IBUFFX4_RVT U1448 ( .A(n506), .Y(n504) );
  IBUFFX4_RVT U1449 ( .A(n505), .Y(n506) );
  INVX1_RVT U1450 ( .A(net30010), .Y(\u_div/PartRem[26][3] ) );
  MUX21X1_RVT U1451 ( .A1(net29991), .A2(net31079), .S0(n145), .Y(net30010) );
  INVX1_RVT U1452 ( .A(net30011), .Y(\u_div/PartRem[26][2] ) );
  MUX21X1_RVT U1453 ( .A1(net29993), .A2(net31099), .S0(n143), .Y(net30011) );
  INVX1_RVT U1454 ( .A(net30014), .Y(\u_div/PartRem[26][1] ) );
  MUX21X1_RVT U1455 ( .A1(net31738), .A2(net37253), .S0(n151), .Y(net30014) );
  OR2X1_RVT U1456 ( .A1(net32406), .A2(a[25]), .Y(\u_div/CryTmp[25][1] ) );
  INVX1_RVT U1457 ( .A(net30005), .Y(\u_div/PartRem[26][8] ) );
  MUX21X1_RVT U1458 ( .A1(net29986), .A2(net30962), .S0(n143), .Y(net30005) );
  OR2X2_RVT U1459 ( .A1(net31315), .A2(n502), .Y(net31317) );
  OR2X1_RVT U1460 ( .A1(net31814), .A2(net31844), .Y(net31315) );
  IBUFFX16_RVT U1461 ( .A(\u_div/CryTmp[25][22] ), .Y(n502) );
  INVX0_RVT U1462 ( .A(net30012), .Y(\u_div/PartRem[26][21] ) );
  MUX21X1_RVT U1463 ( .A1(net29992), .A2(net30080), .S0(n144), .Y(net30012) );
  INVX1_RVT U1464 ( .A(net31872), .Y(net31856) );
  IBUFFX16_RVT U1465 ( .A(net30013), .Y(\u_div/PartRem[26][20] ) );
  MUX21X1_RVT U1466 ( .A1(net29994), .A2(net30143), .S0(n148), .Y(net30013) );
  INVX1_RVT U1467 ( .A(net31896), .Y(net31884) );
  MUX21X1_RVT U1468 ( .A1(net29995), .A2(net30203), .S0(n143), .Y(net30015) );
  MUX21X1_RVT U1469 ( .A1(net29996), .A2(net30251), .S0(n153), .Y(net30016) );
  NBUFFX8_RVT U1470 ( .A(\u_div/CryTmp[25][18] ), .Y(n517) );
  MUX21X1_RVT U1471 ( .A1(net29997), .A2(net30494), .S0(quotient[26]), .Y(
        net30017) );
  INVX1_RVT U1472 ( .A(net30018), .Y(\u_div/PartRem[26][16] ) );
  MUX21X1_RVT U1473 ( .A1(net29998), .A2(net30542), .S0(n149), .Y(net30018) );
  INVX1_RVT U1474 ( .A(net30019), .Y(\u_div/PartRem[26][15] ) );
  MUX21X1_RVT U1475 ( .A1(net29999), .A2(net30590), .S0(n144), .Y(net30019) );
  IBUFFX4_RVT U1476 ( .A(net30020), .Y(\u_div/PartRem[26][14] ) );
  MUX21X1_RVT U1477 ( .A1(net30000), .A2(net30638), .S0(n152), .Y(net30020) );
  INVX0_RVT U1478 ( .A(\u_div/SumTmp[25][20] ), .Y(net30142) );
  INVX0_RVT U1479 ( .A(\u_div/SumTmp[25][19] ), .Y(net30202) );
  INVX0_RVT U1480 ( .A(\u_div/SumTmp[25][18] ), .Y(net30250) );
  INVX0_RVT U1481 ( .A(\u_div/SumTmp[25][17] ), .Y(net30493) );
  INVX0_RVT U1482 ( .A(\u_div/SumTmp[25][16] ), .Y(net30541) );
  INVX0_RVT U1483 ( .A(\u_div/SumTmp[25][15] ), .Y(net30589) );
  IBUFFX16_RVT U1484 ( .A(\u_div/SumTmp[25][14] ), .Y(net30637) );
  INVX1_RVT U1485 ( .A(\u_div/SumTmp[25][11] ), .Y(net30781) );
  INVX1_RVT U1486 ( .A(\u_div/SumTmp[25][10] ), .Y(net30829) );
  INVX1_RVT U1487 ( .A(\u_div/SumTmp[26][8] ), .Y(net30878) );
  MUX21X1_RVT U1488 ( .A1(n549), .A2(net30776), .S0(net32598), .Y(n556) );
  IBUFFX4_RVT U1489 ( .A(\u_div/PartRem[20][16] ), .Y(n589) );
  MUX21X1_RVT U1490 ( .A1(n550), .A2(net30824), .S0(net32598), .Y(net30277) );
  INVX4_RVT U1491 ( .A(n585), .Y(n586) );
  IBUFFX4_RVT U1492 ( .A(\u_div/PartRem[20][15] ), .Y(n585) );
  INVX1_RVT U1493 ( .A(net30278), .Y(\u_div/PartRem[20][15] ) );
  MUX21X1_RVT U1494 ( .A1(n551), .A2(net30872), .S0(net32598), .Y(net30278) );
  INVX1_RVT U1495 ( .A(net32024), .Y(net32014) );
  INVX4_RVT U1496 ( .A(n587), .Y(n588) );
  MUX21X1_RVT U1497 ( .A1(n552), .A2(net30956), .S0(net46961), .Y(net30279) );
  INVX1_RVT U1498 ( .A(b[14]), .Y(net32044) );
  IBUFFX16_RVT U1499 ( .A(\u_div/CryTmp[19][14] ), .Y(n568) );
  INVX1_RVT U1500 ( .A(net30280), .Y(\u_div/PartRem[20][13] ) );
  MUX21X1_RVT U1501 ( .A1(n553), .A2(net30982), .S0(net44969), .Y(net30280) );
  INVX1_RVT U1502 ( .A(net32076), .Y(net32066) );
  INVX1_RVT U1503 ( .A(net30281), .Y(\u_div/PartRem[20][12] ) );
  MUX21X1_RVT U1504 ( .A1(n554), .A2(net31006), .S0(net44969), .Y(net30281) );
  INVX1_RVT U1505 ( .A(net32104), .Y(net32090) );
  INVX1_RVT U1506 ( .A(net30282), .Y(\u_div/PartRem[20][11] ) );
  MUX21X1_RVT U1507 ( .A1(n555), .A2(net31029), .S0(net44969), .Y(net30282) );
  INVX1_RVT U1508 ( .A(net32128), .Y(net32116) );
  MUX21X1_RVT U1509 ( .A1(n540), .A2(net31051), .S0(net44969), .Y(net30283) );
  IBUFFX16_RVT U1510 ( .A(\u_div/CryTmp[19][10] ), .Y(n563) );
  INVX1_RVT U1511 ( .A(net30237), .Y(\u_div/PartRem[20][9] ) );
  INVX1_RVT U1512 ( .A(net30238), .Y(\u_div/PartRem[20][8] ) );
  MUX21X1_RVT U1513 ( .A1(n542), .A2(net31093), .S0(net44969), .Y(net30238) );
  INVX1_RVT U1514 ( .A(net30239), .Y(\u_div/PartRem[20][7] ) );
  MUX21X1_RVT U1515 ( .A1(n543), .A2(net31112), .S0(net44969), .Y(net30239) );
  INVX1_RVT U1516 ( .A(net30240), .Y(\u_div/PartRem[20][6] ) );
  MUX21X1_RVT U1517 ( .A1(n544), .A2(net31130), .S0(net44969), .Y(net30240) );
  INVX1_RVT U1518 ( .A(net32264), .Y(net32252) );
  INVX1_RVT U1519 ( .A(net30241), .Y(\u_div/PartRem[20][5] ) );
  MUX21X1_RVT U1520 ( .A1(n545), .A2(net31147), .S0(net44969), .Y(net30241) );
  INVX1_RVT U1521 ( .A(net32300), .Y(net32282) );
  INVX1_RVT U1522 ( .A(net30242), .Y(\u_div/PartRem[20][4] ) );
  MUX21X1_RVT U1523 ( .A1(n546), .A2(net31163), .S0(net44969), .Y(net30242) );
  INVX1_RVT U1524 ( .A(net32324), .Y(net32312) );
  INVX1_RVT U1525 ( .A(net30243), .Y(\u_div/PartRem[20][3] ) );
  MUX21X1_RVT U1526 ( .A1(n547), .A2(net31178), .S0(net44969), .Y(net30243) );
  INVX1_RVT U1527 ( .A(net32352), .Y(net32336) );
  INVX1_RVT U1528 ( .A(net30244), .Y(\u_div/PartRem[20][2] ) );
  MUX21X1_RVT U1529 ( .A1(n548), .A2(net31191), .S0(net44969), .Y(net30244) );
  INVX1_RVT U1530 ( .A(b[2]), .Y(net32364) );
  INVX1_RVT U1531 ( .A(b[1]), .Y(net32384) );
  INVX1_RVT U1532 ( .A(net30273), .Y(\u_div/PartRem[20][1] ) );
  NAND2X0_RVT U1533 ( .A1(net44969), .A2(\*cell*33669/net34055 ), .Y(net30273)
         );
  INVX1_RVT U1534 ( .A(b[0]), .Y(\u_div/CryTmp[22][1] ) );
  INVX0_RVT U1535 ( .A(\u_div/SumTmp[19][17] ), .Y(net30775) );
  INVX0_RVT U1536 ( .A(\u_div/SumTmp[20][16] ), .Y(net30776) );
  INVX1_RVT U1537 ( .A(n549), .Y(\u_div/PartRem[21][16] ) );
  MUX21X1_RVT U1538 ( .A1(net30185), .A2(net30825), .S0(n209), .Y(n550) );
  MUX21X1_RVT U1539 ( .A1(net30186), .A2(net30873), .S0(n205), .Y(n551) );
  MUX21X1_RVT U1540 ( .A1(net30187), .A2(net30957), .S0(n204), .Y(n552) );
  MUX21X1_RVT U1541 ( .A1(net30189), .A2(net31007), .S0(n200), .Y(n554) );
  INVX1_RVT U1542 ( .A(n555), .Y(\u_div/PartRem[21][10] ) );
  MUX21X1_RVT U1543 ( .A1(net30131), .A2(net31030), .S0(n202), .Y(n555) );
  INVX2_RVT U1544 ( .A(n580), .Y(n581) );
  IBUFFX4_RVT U1545 ( .A(\u_div/CryTmp[20][8] ), .Y(n580) );
  INVX1_RVT U1546 ( .A(n542), .Y(\u_div/PartRem[21][7] ) );
  MUX21X1_RVT U1547 ( .A1(net30134), .A2(net31094), .S0(n203), .Y(n542) );
  IBUFFX16_RVT U1548 ( .A(n543), .Y(\u_div/PartRem[21][6] ) );
  MUX21X1_RVT U1549 ( .A1(net30135), .A2(net31113), .S0(n204), .Y(n543) );
  INVX1_RVT U1550 ( .A(n544), .Y(\u_div/PartRem[21][5] ) );
  MUX21X1_RVT U1551 ( .A1(net30136), .A2(net31131), .S0(n202), .Y(n544) );
  INVX1_RVT U1552 ( .A(n545), .Y(\u_div/PartRem[21][4] ) );
  MUX21X1_RVT U1553 ( .A1(net30137), .A2(net31148), .S0(n201), .Y(n545) );
  INVX1_RVT U1554 ( .A(n546), .Y(\u_div/PartRem[21][3] ) );
  MUX21X1_RVT U1555 ( .A1(net30138), .A2(net31164), .S0(n200), .Y(n546) );
  INVX1_RVT U1556 ( .A(n547), .Y(\u_div/PartRem[21][2] ) );
  MUX21X1_RVT U1557 ( .A1(net30179), .A2(net31179), .S0(n203), .Y(n547) );
  INVX1_RVT U1558 ( .A(n548), .Y(n565) );
  NAND2X0_RVT U1559 ( .A1(n199), .A2(\*cell*33672/net34065 ), .Y(n548) );
  MUX21X1_RVT U1560 ( .A1(n556), .A2(net30775), .S0(net32592), .Y(net30517) );
  INVX0_RVT U1561 ( .A(\u_div/SumTmp[20][15] ), .Y(net30824) );
  INVX0_RVT U1562 ( .A(\u_div/SumTmp[20][13] ), .Y(net30956) );
  INVX0_RVT U1563 ( .A(\u_div/SumTmp[20][12] ), .Y(net30982) );
  MUX21X1_RVT U1564 ( .A1(net30130), .A2(net30984), .S0(net32608), .Y(net30188) );
  INVX0_RVT U1565 ( .A(\u_div/SumTmp[21][11] ), .Y(net30983) );
  INVX1_RVT U1566 ( .A(net30188), .Y(\u_div/PartRem[22][11] ) );
  INVX1_RVT U1567 ( .A(net30189), .Y(\u_div/PartRem[22][10] ) );
  MUX21X1_RVT U1568 ( .A1(net30069), .A2(net31008), .S0(net32608), .Y(net30189) );
  MUX21X1_RVT U1569 ( .A1(net30070), .A2(net31031), .S0(net32608), .Y(net30131) );
  MUX21X1_RVT U1570 ( .A1(net30071), .A2(net31053), .S0(net32608), .Y(net30132) );
  MUX21X1_RVT U1571 ( .A1(net30072), .A2(net31075), .S0(net32608), .Y(net30133) );
  INVX1_RVT U1572 ( .A(net30134), .Y(\u_div/PartRem[22][6] ) );
  INVX4_RVT U1573 ( .A(n561), .Y(n562) );
  IBUFFX16_RVT U1574 ( .A(\u_div/CryTmp[21][5] ), .Y(n561) );
  INVX1_RVT U1575 ( .A(net30136), .Y(\u_div/PartRem[22][4] ) );
  MUX21X1_RVT U1576 ( .A1(n534), .A2(net31132), .S0(net32608), .Y(net30136) );
  INVX1_RVT U1577 ( .A(net30137), .Y(\u_div/PartRem[22][3] ) );
  MUX21X1_RVT U1578 ( .A1(n535), .A2(net31149), .S0(net32608), .Y(net30137) );
  INVX1_RVT U1579 ( .A(net30138), .Y(\u_div/PartRem[22][2] ) );
  MUX21X1_RVT U1580 ( .A1(n536), .A2(net31165), .S0(net32608), .Y(net30138) );
  INVX1_RVT U1581 ( .A(net30179), .Y(\u_div/PartRem[22][1] ) );
  NAND2X0_RVT U1582 ( .A1(net32608), .A2(\*cell*33675/net34075 ), .Y(net30179)
         );
  MUX21X1_RVT U1583 ( .A1(\u_div/SumTmp[22][4] ), .A2(\u_div/PartRem[23][4] ), 
        .S0(n560), .Y(net46688) );
  IBUFFX16_RVT U1584 ( .A(\u_div/CryTmp[21][12] ), .Y(net49112) );
  INVX0_RVT U1585 ( .A(\u_div/SumTmp[21][10] ), .Y(net31007) );
  INVX0_RVT U1586 ( .A(\u_div/SumTmp[21][9] ), .Y(net31030) );
  INVX0_RVT U1587 ( .A(\u_div/SumTmp[21][8] ), .Y(net31052) );
  INVX0_RVT U1588 ( .A(\u_div/SumTmp[21][7] ), .Y(net31074) );
  MUX21X1_RVT U1589 ( .A1(n523), .A2(net31096), .S0(quotient[23]), .Y(n533) );
  INVX0_RVT U1590 ( .A(\u_div/SumTmp[22][5] ), .Y(n557) );
  INVX2_RVT U1591 ( .A(net30074), .Y(\u_div/PartRem[23][4] ) );
  MUX21X1_RVT U1592 ( .A1(n524), .A2(net31133), .S0(quotient[23]), .Y(n534) );
  MUX21X1_RVT U1593 ( .A1(n528), .A2(net31150), .S0(quotient[23]), .Y(n535) );
  INVX1_RVT U1594 ( .A(n536), .Y(\u_div/PartRem[23][1] ) );
  MUX21X2_RVT U1595 ( .A1(net31786), .A2(net37228), .S0(quotient[23]), .Y(n536) );
  INVX1_RVT U1596 ( .A(n560), .Y(net32608) );
  NOR2X0_RVT U1597 ( .A1(\u_div/CryTmp[22][24] ), .A2(\u_div/PartRem[23][24] ), 
        .Y(n560) );
  INVX1_RVT U1598 ( .A(n537), .Y(\u_div/PartRem[23][23] ) );
  IBUFFX32_RVT U1599 ( .A(\u_div/CryTmp[22][23] ), .Y(n576) );
  MUX21X1_RVT U1600 ( .A1(n526), .A2(net30200), .S0(quotient[23]), .Y(net30117) );
  INVX1_RVT U1601 ( .A(net31844), .Y(net31828) );
  IBUFFX16_RVT U1602 ( .A(net30118), .Y(\u_div/PartRem[23][21] ) );
  MUX21X1_RVT U1603 ( .A1(n527), .A2(net30248), .S0(n1240), .Y(net30118) );
  IBUFFX16_RVT U1604 ( .A(net30119), .Y(\u_div/PartRem[23][20] ) );
  MUX21X1_RVT U1605 ( .A1(n529), .A2(net30491), .S0(n1240), .Y(net30119) );
  IBUFFX16_RVT U1606 ( .A(net30121), .Y(\u_div/PartRem[23][19] ) );
  MUX21X1_RVT U1607 ( .A1(n530), .A2(net30539), .S0(n1240), .Y(net30121) );
  INVX1_RVT U1608 ( .A(net31922), .Y(net31912) );
  IBUFFX16_RVT U1609 ( .A(net30122), .Y(\u_div/PartRem[23][18] ) );
  MUX21X1_RVT U1610 ( .A1(n531), .A2(net30587), .S0(quotient[23]), .Y(net30122) );
  IBUFFX4_RVT U1611 ( .A(n578), .Y(n579) );
  IBUFFX32_RVT U1612 ( .A(\u_div/CryTmp[22][18] ), .Y(n578) );
  MUX21X1_RVT U1613 ( .A1(n532), .A2(net30635), .S0(quotient[23]), .Y(net30123) );
  NAND3X0_RVT U1614 ( .A1(n582), .A2(n583), .A3(n584), .Y(
        \u_div/CryTmp[22][17] ) );
  NAND2X0_RVT U1615 ( .A1(n33), .A2(net31982), .Y(n582) );
  NAND3X0_RVT U1616 ( .A1(net49309), .A2(net49310), .A3(net49311), .Y(
        \u_div/CryTmp[22][16] ) );
  NAND2X0_RVT U1617 ( .A1(net31982), .A2(\u_div/CryTmp[22][16] ), .Y(n584) );
  INVX1_RVT U1618 ( .A(net31814), .Y(net31802) );
  MUX21X1_RVT U1619 ( .A1(n559), .A2(\u_div/SumTmp[23][23] ), .S0(quotient[23]), .Y(\u_div/PartRem[23][24] ) );
  INVX1_RVT U1620 ( .A(n525), .Y(\u_div/PartRem[24][22] ) );
  MUX21X1_RVT U1621 ( .A1(n522), .A2(n539), .S0(net47709), .Y(n525) );
  MUX21X1_RVT U1622 ( .A1(net30035), .A2(net30201), .S0(net47709), .Y(n526) );
  IBUFFX16_RVT U1623 ( .A(n527), .Y(\u_div/PartRem[24][20] ) );
  MUX21X1_RVT U1624 ( .A1(net30037), .A2(net30249), .S0(net32620), .Y(n527) );
  IBUFFX16_RVT U1625 ( .A(n529), .Y(\u_div/PartRem[24][19] ) );
  MUX21X1_RVT U1626 ( .A1(net30038), .A2(net30492), .S0(net32620), .Y(n529) );
  IBUFFX16_RVT U1627 ( .A(n530), .Y(\u_div/PartRem[24][18] ) );
  IBUFFX16_RVT U1628 ( .A(n531), .Y(\u_div/PartRem[24][17] ) );
  IBUFFX16_RVT U1629 ( .A(net30064), .Y(\u_div/PartRem[24][14] ) );
  INVX1_RVT U1630 ( .A(net30065), .Y(\u_div/PartRem[24][13] ) );
  MUX21X1_RVT U1631 ( .A1(net30044), .A2(net30780), .S0(net32620), .Y(net30065) );
  INVX1_RVT U1632 ( .A(net30066), .Y(\u_div/PartRem[24][12] ) );
  MUX21X1_RVT U1633 ( .A1(net30045), .A2(net30828), .S0(net32620), .Y(net30066) );
  INVX1_RVT U1634 ( .A(net30067), .Y(\u_div/PartRem[24][11] ) );
  MUX21X1_RVT U1635 ( .A1(net41435), .A2(net30876), .S0(net47709), .Y(net30067) );
  INVX1_RVT U1636 ( .A(net30068), .Y(\u_div/PartRem[24][10] ) );
  MUX21X1_RVT U1637 ( .A1(net30025), .A2(net30960), .S0(net32620), .Y(net30068) );
  INVX1_RVT U1638 ( .A(net30047), .Y(\u_div/PartRem[24][9] ) );
  MUX21X1_RVT U1639 ( .A1(net30026), .A2(net30986), .S0(net32620), .Y(net30047) );
  INVX1_RVT U1640 ( .A(net30048), .Y(\u_div/PartRem[24][8] ) );
  MUX21X1_RVT U1641 ( .A1(net30027), .A2(net31010), .S0(net32620), .Y(net30048) );
  INVX1_RVT U1642 ( .A(net30049), .Y(\u_div/PartRem[24][7] ) );
  MUX21X1_RVT U1643 ( .A1(net30028), .A2(net31033), .S0(net47709), .Y(net30049) );
  INVX1_RVT U1644 ( .A(net30050), .Y(\u_div/PartRem[24][6] ) );
  MUX21X1_RVT U1645 ( .A1(net30029), .A2(net31055), .S0(net47709), .Y(net30050) );
  INVX1_RVT U1646 ( .A(net30051), .Y(\u_div/PartRem[24][5] ) );
  MUX21X1_RVT U1647 ( .A1(net30030), .A2(net31077), .S0(net47709), .Y(net30051) );
  INVX1_RVT U1648 ( .A(n523), .Y(\u_div/PartRem[24][4] ) );
  MUX21X1_RVT U1649 ( .A1(net30031), .A2(net31097), .S0(net47709), .Y(n523) );
  INVX1_RVT U1650 ( .A(net30053), .Y(\u_div/PartRem[24][3] ) );
  MUX21X1_RVT U1651 ( .A1(net30032), .A2(net31116), .S0(net47709), .Y(net30053) );
  INVX1_RVT U1652 ( .A(n524), .Y(\u_div/PartRem[24][2] ) );
  MUX21X1_RVT U1653 ( .A1(net30036), .A2(net31134), .S0(net47709), .Y(n524) );
  INVX1_RVT U1654 ( .A(n528), .Y(\u_div/PartRem[24][1] ) );
  MUX21X1_RVT U1655 ( .A1(net31770), .A2(net37229), .S0(net47709), .Y(n528) );
  OR2X1_RVT U1656 ( .A1(\u_div/CryTmp[22][1] ), .A2(a[23]), .Y(
        \u_div/CryTmp[23][1] ) );
  IBUFFX16_RVT U1657 ( .A(n1240), .Y(n558) );
  IBUFFX16_RVT U1658 ( .A(\u_div/SumTmp[23][22] ), .Y(n538) );
  MUX21X1_RVT U1659 ( .A1(net30013), .A2(net30142), .S0(quotient[25]), .Y(n522) );
  INVX0_RVT U1660 ( .A(\u_div/SumTmp[24][21] ), .Y(n539) );
  INVX1_RVT U1661 ( .A(n522), .Y(\u_div/PartRem[25][21] ) );
  INVX1_RVT U1662 ( .A(net31872), .Y(net31854) );
  IBUFFX16_RVT U1663 ( .A(net30035), .Y(\u_div/PartRem[25][20] ) );
  MUX21X1_RVT U1664 ( .A1(net30015), .A2(net30202), .S0(quotient[25]), .Y(
        net30035) );
  MUX21X1_RVT U1665 ( .A1(n525), .A2(n538), .S0(quotient[23]), .Y(n537) );
  INVX0_RVT U1666 ( .A(\u_div/SumTmp[24][20] ), .Y(net30201) );
  INVX1_RVT U1667 ( .A(n617), .Y(\u_div/PartRem[17][1] ) );
  NAND2X0_RVT U1668 ( .A1(n158), .A2(\*cell*33699/net34155 ), .Y(n617) );
  INVX0_RVT U1669 ( .A(net30918), .Y(\*cell*33699/net34155 ) );
  INVX0_RVT U1670 ( .A(\u_div/SumTmp[17][0] ), .Y(net30918) );
  INVX0_RVT U1671 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[17][0] ) );
  MUX21X1_RVT U1672 ( .A1(n617), .A2(net30917), .S0(n11), .Y(net30627) );
  NOR2X2_RVT U1673 ( .A1(\u_div/PartRem[18][24] ), .A2(\u_div/CryTmp[17][24] ), 
        .Y(net38346) );
  MUX21X1_RVT U1674 ( .A1(\u_div/PartRem[19][23] ), .A2(\u_div/SumTmp[18][23] ), .S0(n636), .Y(\u_div/PartRem[18][24] ) );
  INVX1_RVT U1675 ( .A(net30534), .Y(\u_div/PartRem[19][23] ) );
  INVX2_RVT U1676 ( .A(net30512), .Y(\u_div/PartRem[19][22] ) );
  INVX1_RVT U1677 ( .A(n605), .Y(\u_div/PartRem[19][21] ) );
  MUX21X1_RVT U1678 ( .A1(n595), .A2(n619), .S0(net32590), .Y(n605) );
  INVX1_RVT U1679 ( .A(n606), .Y(\u_div/PartRem[19][20] ) );
  MUX21X1_RVT U1680 ( .A1(n596), .A2(n621), .S0(net32592), .Y(n606) );
  INVX1_RVT U1681 ( .A(n608), .Y(\u_div/PartRem[19][19] ) );
  MUX21X1_RVT U1682 ( .A1(net30275), .A2(net30727), .S0(net32592), .Y(n608) );
  INVX1_RVT U1683 ( .A(net30517), .Y(\u_div/PartRem[19][18] ) );
  INVX1_RVT U1684 ( .A(n610), .Y(\u_div/PartRem[19][16] ) );
  MUX21X1_RVT U1685 ( .A1(net30278), .A2(net30871), .S0(net32590), .Y(n610) );
  INVX1_RVT U1686 ( .A(net31998), .Y(net31984) );
  INVX1_RVT U1687 ( .A(n611), .Y(\u_div/PartRem[19][15] ) );
  IBUFFX16_RVT U1688 ( .A(\u_div/CryTmp[18][15] ), .Y(n625) );
  INVX1_RVT U1689 ( .A(n612), .Y(\u_div/PartRem[19][14] ) );
  MUX21X1_RVT U1690 ( .A1(net30280), .A2(net30981), .S0(net32590), .Y(n612) );
  INVX1_RVT U1691 ( .A(n613), .Y(\u_div/PartRem[19][13] ) );
  MUX21X1_RVT U1692 ( .A1(net30281), .A2(net31005), .S0(net32590), .Y(n613) );
  INVX1_RVT U1693 ( .A(n614), .Y(\u_div/PartRem[19][12] ) );
  MUX21X1_RVT U1694 ( .A1(net30282), .A2(net31028), .S0(net32590), .Y(n614) );
  INVX1_RVT U1695 ( .A(n615), .Y(\u_div/PartRem[19][11] ) );
  MUX21X1_RVT U1696 ( .A1(net30283), .A2(net31050), .S0(net32590), .Y(n615) );
  INVX1_RVT U1697 ( .A(n616), .Y(\u_div/PartRem[19][10] ) );
  MUX21X1_RVT U1698 ( .A1(net30237), .A2(net31072), .S0(net32590), .Y(n616) );
  INVX1_RVT U1699 ( .A(n597), .Y(\u_div/PartRem[19][9] ) );
  MUX21X1_RVT U1700 ( .A1(net30238), .A2(net31092), .S0(net32590), .Y(n597) );
  INVX1_RVT U1701 ( .A(n598), .Y(\u_div/PartRem[19][8] ) );
  MUX21X1_RVT U1702 ( .A1(net30239), .A2(net31111), .S0(net32590), .Y(n598) );
  INVX1_RVT U1703 ( .A(n599), .Y(\u_div/PartRem[19][7] ) );
  MUX21X1_RVT U1704 ( .A1(net30240), .A2(net31129), .S0(net32590), .Y(n599) );
  INVX1_RVT U1705 ( .A(n600), .Y(\u_div/PartRem[19][6] ) );
  MUX21X1_RVT U1706 ( .A1(net30241), .A2(net31146), .S0(net32590), .Y(n600) );
  INVX1_RVT U1707 ( .A(n601), .Y(\u_div/PartRem[19][5] ) );
  MUX21X1_RVT U1708 ( .A1(net30242), .A2(net31162), .S0(net32592), .Y(n601) );
  INVX1_RVT U1709 ( .A(n602), .Y(\u_div/PartRem[19][4] ) );
  MUX21X1_RVT U1710 ( .A1(net30243), .A2(net31177), .S0(net32592), .Y(n602) );
  INVX1_RVT U1711 ( .A(n603), .Y(\u_div/PartRem[19][3] ) );
  MUX21X1_RVT U1712 ( .A1(net30244), .A2(net31190), .S0(n212), .Y(n603) );
  MUX21X1_RVT U1713 ( .A1(net30273), .A2(net31202), .S0(n211), .Y(n604) );
  INVX1_RVT U1714 ( .A(n607), .Y(\u_div/PartRem[19][1] ) );
  NAND2X0_RVT U1715 ( .A1(n211), .A2(\*cell*33666/net34045 ), .Y(n607) );
  INVX1_RVT U1716 ( .A(net45669), .Y(n636) );
  INVX1_RVT U1717 ( .A(net30560), .Y(\u_div/PartRem[18][21] ) );
  MUX21X1_RVT U1718 ( .A1(n606), .A2(n620), .S0(net45665), .Y(net30560) );
  IBUFFX4_RVT U1719 ( .A(n641), .Y(n642) );
  INVX1_RVT U1720 ( .A(\u_div/CryTmp[17][20] ), .Y(n641) );
  INVX1_RVT U1721 ( .A(net30563), .Y(\u_div/PartRem[18][19] ) );
  MUX21X1_RVT U1722 ( .A1(net30517), .A2(n623), .S0(net45671), .Y(net30563) );
  IBUFFX16_RVT U1723 ( .A(\u_div/CryTmp[17][19] ), .Y(n631) );
  INVX1_RVT U1724 ( .A(net30564), .Y(\u_div/PartRem[18][18] ) );
  MUX21X1_RVT U1725 ( .A1(n609), .A2(n624), .S0(n637), .Y(net30564) );
  INVX1_RVT U1726 ( .A(net30565), .Y(\u_div/PartRem[18][17] ) );
  MUX21X1_RVT U1727 ( .A1(n610), .A2(net30870), .S0(net45677), .Y(net30565) );
  INVX1_RVT U1728 ( .A(net31972), .Y(net31962) );
  INVX1_RVT U1729 ( .A(net30566), .Y(\u_div/PartRem[18][16] ) );
  MUX21X1_RVT U1730 ( .A1(n611), .A2(net30954), .S0(net45677), .Y(net30566) );
  IBUFFX16_RVT U1731 ( .A(net30567), .Y(\u_div/PartRem[18][15] ) );
  MUX21X1_RVT U1732 ( .A1(n612), .A2(net30980), .S0(n635), .Y(net30567) );
  IBUFFX16_RVT U1733 ( .A(net30568), .Y(\u_div/PartRem[18][14] ) );
  MUX21X1_RVT U1734 ( .A1(n613), .A2(net31004), .S0(net45678), .Y(net30568) );
  IBUFFX16_RVT U1735 ( .A(\u_div/CryTmp[17][14] ), .Y(n629) );
  INVX1_RVT U1736 ( .A(net30569), .Y(\u_div/PartRem[18][13] ) );
  MUX21X1_RVT U1737 ( .A1(n614), .A2(net31027), .S0(n637), .Y(net30569) );
  INVX1_RVT U1738 ( .A(net30570), .Y(\u_div/PartRem[18][12] ) );
  MUX21X1_RVT U1739 ( .A1(n615), .A2(net31049), .S0(n635), .Y(net30570) );
  INVX1_RVT U1740 ( .A(net30571), .Y(\u_div/PartRem[18][11] ) );
  MUX21X1_RVT U1741 ( .A1(n616), .A2(net31071), .S0(net45665), .Y(net30571) );
  IBUFFX16_RVT U1742 ( .A(net30572), .Y(\u_div/PartRem[18][10] ) );
  MUX21X1_RVT U1743 ( .A1(n597), .A2(net31091), .S0(net45678), .Y(net30572) );
  IBUFFX16_RVT U1744 ( .A(net30526), .Y(\u_div/PartRem[18][9] ) );
  MUX21X1_RVT U1745 ( .A1(n598), .A2(net31110), .S0(net45677), .Y(net30526) );
  IBUFFX16_RVT U1746 ( .A(net30527), .Y(\u_div/PartRem[18][8] ) );
  MUX21X1_RVT U1747 ( .A1(n599), .A2(net31128), .S0(n636), .Y(net30527) );
  IBUFFX4_RVT U1748 ( .A(n639), .Y(n640) );
  IBUFFX2_RVT U1749 ( .A(\u_div/CryTmp[17][8] ), .Y(n639) );
  INVX4_RVT U1750 ( .A(n627), .Y(n628) );
  IBUFFX16_RVT U1751 ( .A(\u_div/CryTmp[17][7] ), .Y(n627) );
  INVX1_RVT U1752 ( .A(net30529), .Y(\u_div/PartRem[18][6] ) );
  MUX21X1_RVT U1753 ( .A1(n601), .A2(net31161), .S0(n635), .Y(net30529) );
  INVX1_RVT U1754 ( .A(net30530), .Y(\u_div/PartRem[18][5] ) );
  MUX21X1_RVT U1755 ( .A1(n602), .A2(net31176), .S0(n636), .Y(net30530) );
  INVX1_RVT U1756 ( .A(net30531), .Y(\u_div/PartRem[18][4] ) );
  MUX21X1_RVT U1757 ( .A1(n603), .A2(net31189), .S0(net45671), .Y(net30531) );
  INVX1_RVT U1758 ( .A(net30532), .Y(\u_div/PartRem[18][3] ) );
  MUX21X1_RVT U1759 ( .A1(n604), .A2(net31201), .S0(n635), .Y(net30532) );
  INVX1_RVT U1760 ( .A(net30533), .Y(\u_div/PartRem[18][2] ) );
  INVX1_RVT U1761 ( .A(net30562), .Y(\u_div/PartRem[18][1] ) );
  NAND2X0_RVT U1762 ( .A1(net45671), .A2(\*cell*33702/net34165 ), .Y(net30562)
         );
  INVX2_RVT U1763 ( .A(net30561), .Y(\u_div/PartRem[18][20] ) );
  MUX21X2_RVT U1764 ( .A1(n608), .A2(n622), .S0(n637), .Y(net30561) );
  INVX2_RVT U1765 ( .A(net30559), .Y(\u_div/PartRem[18][22] ) );
  MUX21X2_RVT U1766 ( .A1(n605), .A2(n618), .S0(net45665), .Y(net30559) );
  INVX4_RVT U1767 ( .A(net38346), .Y(net32580) );
  MUX21X1_RVT U1768 ( .A1(n638), .A2(\u_div/SumTmp[17][23] ), .S0(n158), .Y(
        \u_div/PartRem[17][24] ) );
  INVX0_RVT U1769 ( .A(\u_div/SumTmp[17][22] ), .Y(net30629) );
  INVX0_RVT U1770 ( .A(\u_div/SumTmp[17][21] ), .Y(net30677) );
  INVX0_RVT U1771 ( .A(\u_div/SumTmp[17][20] ), .Y(net30725) );
  INVX0_RVT U1772 ( .A(\u_div/SumTmp[18][19] ), .Y(n622) );
  INVX1_RVT U1773 ( .A(net45669), .Y(n637) );
  MUX21X1_RVT U1774 ( .A1(net30561), .A2(net30725), .S0(n157), .Y(net30607) );
  MUX21X1_RVT U1775 ( .A1(\u_div/PartRem[20][23] ), .A2(\u_div/SumTmp[19][23] ), .S0(net32590), .Y(\u_div/PartRem[19][24] ) );
  INVX0_RVT U1776 ( .A(\u_div/SumTmp[18][21] ), .Y(n618) );
  INVX0_RVT U1777 ( .A(\u_div/SumTmp[18][20] ), .Y(n620) );
  INVX0_RVT U1778 ( .A(\u_div/SumTmp[18][18] ), .Y(n623) );
  INVX0_RVT U1779 ( .A(\u_div/SumTmp[18][17] ), .Y(n624) );
  INVX0_RVT U1780 ( .A(\u_div/SumTmp[19][16] ), .Y(net30823) );
  INVX0_RVT U1781 ( .A(net38344), .Y(net32592) );
  INVX1_RVT U1782 ( .A(net30487), .Y(\u_div/PartRem[20][23] ) );
  INVX1_RVT U1783 ( .A(net30270), .Y(\u_div/PartRem[20][22] ) );
  MUX21X1_RVT U1784 ( .A1(n591), .A2(net30536), .S0(net32598), .Y(net30270) );
  INVX1_RVT U1785 ( .A(net30271), .Y(\u_div/PartRem[20][21] ) );
  MUX21X1_RVT U1786 ( .A1(n592), .A2(net30584), .S0(net32598), .Y(net30271) );
  INVX1_RVT U1787 ( .A(n595), .Y(\u_div/PartRem[20][20] ) );
  INVX1_RVT U1788 ( .A(n596), .Y(\u_div/PartRem[20][19] ) );
  MUX21X1_RVT U1789 ( .A1(n594), .A2(net30680), .S0(net32598), .Y(n596) );
  INVX1_RVT U1790 ( .A(net30275), .Y(\u_div/PartRem[20][18] ) );
  MUX21X1_RVT U1791 ( .A1(net30229), .A2(net30728), .S0(net32598), .Y(net30275) );
  MUX21X1_RVT U1792 ( .A1(\u_div/PartRem[21][23] ), .A2(\u_div/SumTmp[20][23] ), .S0(net32598), .Y(\u_div/PartRem[20][24] ) );
  INVX1_RVT U1793 ( .A(net30245), .Y(\u_div/PartRem[21][23] ) );
  INVX1_RVT U1794 ( .A(net30223), .Y(\u_div/PartRem[21][22] ) );
  MUX21X1_RVT U1795 ( .A1(net30177), .A2(net30489), .S0(n208), .Y(net30223) );
  IBUFFX16_RVT U1796 ( .A(\u_div/CryTmp[20][22] ), .Y(n643) );
  MUX21X1_RVT U1797 ( .A1(net30178), .A2(net30537), .S0(n199), .Y(n591) );
  INVX1_RVT U1798 ( .A(n592), .Y(\u_div/PartRem[21][20] ) );
  MUX21X1_RVT U1799 ( .A1(net30180), .A2(net30585), .S0(n195), .Y(n592) );
  MUX21X1_RVT U1800 ( .A1(net30181), .A2(net30633), .S0(n210), .Y(n593) );
  INVX1_RVT U1801 ( .A(n594), .Y(\u_div/PartRem[21][18] ) );
  MUX21X1_RVT U1802 ( .A1(net30182), .A2(net30681), .S0(n207), .Y(n594) );
  INVX1_RVT U1803 ( .A(net30229), .Y(\u_div/PartRem[21][17] ) );
  MUX21X1_RVT U1804 ( .A1(net30183), .A2(net30729), .S0(n193), .Y(net30229) );
  INVX0_RVT U1805 ( .A(\u_div/SumTmp[19][22] ), .Y(net30535) );
  INVX0_RVT U1806 ( .A(\u_div/SumTmp[19][21] ), .Y(net30583) );
  INVX0_RVT U1807 ( .A(\u_div/SumTmp[19][20] ), .Y(n619) );
  INVX0_RVT U1808 ( .A(\u_div/SumTmp[19][19] ), .Y(n621) );
  INVX0_RVT U1809 ( .A(\u_div/SumTmp[19][18] ), .Y(net30727) );
  INVX1_RVT U1810 ( .A(n663), .Y(\u_div/PartRem[15][12] ) );
  MUX21X1_RVT U1811 ( .A1(n662), .A2(n668), .S0(n12), .Y(net30665) );
  IBUFFX16_RVT U1812 ( .A(\u_div/SumTmp[15][11] ), .Y(net31107) );
  INVX1_RVT U1813 ( .A(net30665), .Y(\u_div/PartRem[16][11] ) );
  INVX1_RVT U1814 ( .A(net30666), .Y(\u_div/PartRem[16][10] ) );
  MUX21X1_RVT U1815 ( .A1(n645), .A2(n669), .S0(n20), .Y(net30666) );
  INVX1_RVT U1816 ( .A(net30620), .Y(\u_div/PartRem[16][9] ) );
  MUX21X1_RVT U1817 ( .A1(n646), .A2(n670), .S0(n18), .Y(net30620) );
  INVX1_RVT U1818 ( .A(net30621), .Y(\u_div/PartRem[16][8] ) );
  MUX21X1_RVT U1819 ( .A1(n647), .A2(n671), .S0(n15), .Y(net30621) );
  INVX1_RVT U1820 ( .A(net30622), .Y(\u_div/PartRem[16][7] ) );
  MUX21X1_RVT U1821 ( .A1(n648), .A2(n672), .S0(n13), .Y(net30622) );
  INVX1_RVT U1822 ( .A(net30623), .Y(\u_div/PartRem[16][6] ) );
  MUX21X1_RVT U1823 ( .A1(n649), .A2(n673), .S0(n20), .Y(net30623) );
  INVX1_RVT U1824 ( .A(net30625), .Y(\u_div/PartRem[16][4] ) );
  MUX21X1_RVT U1825 ( .A1(n651), .A2(n675), .S0(n17), .Y(net30625) );
  MUX21X1_RVT U1826 ( .A1(n652), .A2(n664), .S0(n12), .Y(net30626) );
  IBUFFX4_RVT U1827 ( .A(net30627), .Y(\u_div/PartRem[16][2] ) );
  INVX1_RVT U1828 ( .A(net30656), .Y(\u_div/PartRem[16][1] ) );
  NAND2X0_RVT U1829 ( .A1(n13), .A2(\*cell*33696/net34145 ), .Y(net30656) );
  INVX1_RVT U1830 ( .A(net30624), .Y(\u_div/PartRem[16][5] ) );
  MUX21X1_RVT U1831 ( .A1(n650), .A2(n674), .S0(n18), .Y(net30624) );
  MUX21X1_RVT U1832 ( .A1(n663), .A2(net31106), .S0(net47718), .Y(net30757) );
  NOR2X2_RVT U1833 ( .A1(\u_div/CryTmp[15][24] ), .A2(\u_div/PartRem[16][24] ), 
        .Y(net38340) );
  MUX21X1_RVT U1834 ( .A1(net30607), .A2(net30724), .S0(n11), .Y(net30653) );
  MUX21X1_RVT U1835 ( .A1(n653), .A2(net30772), .S0(n5), .Y(net30654) );
  IBUFFX4_RVT U1836 ( .A(net30655), .Y(\u_div/PartRem[16][20] ) );
  MUX21X1_RVT U1837 ( .A1(n654), .A2(net30820), .S0(n16), .Y(net30655) );
  MUX21X1_RVT U1838 ( .A1(n655), .A2(net30868), .S0(n6), .Y(net30657) );
  MUX21X1_RVT U1839 ( .A1(n656), .A2(net30952), .S0(n22), .Y(net30658) );
  INVX1_RVT U1840 ( .A(net31950), .Y(net31940) );
  MUX21X1_RVT U1841 ( .A1(net30613), .A2(net30978), .S0(n15), .Y(n678) );
  MUX21X1_RVT U1842 ( .A1(net30567), .A2(net30979), .S0(n158), .Y(net30613) );
  INVX0_RVT U1843 ( .A(\u_div/SumTmp[16][16] ), .Y(net30978) );
  INVX1_RVT U1844 ( .A(net30661), .Y(\u_div/PartRem[16][15] ) );
  MUX21X1_RVT U1845 ( .A1(n658), .A2(net31025), .S0(n7), .Y(net30661) );
  MUX21X1_RVT U1846 ( .A1(n659), .A2(n665), .S0(quotient[16]), .Y(net30662) );
  MUX21X1_RVT U1847 ( .A1(n660), .A2(n666), .S0(n16), .Y(net30663) );
  MUX21X1_RVT U1848 ( .A1(n661), .A2(n667), .S0(n14), .Y(net30664) );
  INVX1_RVT U1849 ( .A(net30660), .Y(\u_div/PartRem[16][16] ) );
  MUX21X1_RVT U1850 ( .A1(n657), .A2(net31002), .S0(n14), .Y(net30660) );
  MUX21X1_RVT U1851 ( .A1(\u_div/PartRem[17][23] ), .A2(\u_div/SumTmp[16][23] ), .S0(n19), .Y(\u_div/PartRem[16][24] ) );
  INVX1_RVT U1852 ( .A(net30606), .Y(\u_div/PartRem[17][22] ) );
  MUX21X1_RVT U1853 ( .A1(net30560), .A2(net30677), .S0(n158), .Y(net30606) );
  IBUFFX4_RVT U1854 ( .A(\u_div/PartRem[17][21] ), .Y(net52401) );
  INVX1_RVT U1855 ( .A(net30607), .Y(\u_div/PartRem[17][21] ) );
  IBUFFX16_RVT U1856 ( .A(\u_div/CryTmp[16][21] ), .Y(n679) );
  INVX1_RVT U1857 ( .A(n653), .Y(\u_div/PartRem[17][20] ) );
  MUX21X1_RVT U1858 ( .A1(net30563), .A2(net30773), .S0(n158), .Y(n653) );
  INVX1_RVT U1859 ( .A(n654), .Y(\u_div/PartRem[17][19] ) );
  MUX21X1_RVT U1860 ( .A1(net30564), .A2(net30821), .S0(n158), .Y(n654) );
  INVX2_RVT U1861 ( .A(n655), .Y(\u_div/PartRem[17][18] ) );
  MUX21X1_RVT U1862 ( .A1(net30565), .A2(net30869), .S0(n158), .Y(n655) );
  IBUFFX16_RVT U1863 ( .A(n656), .Y(\u_div/PartRem[17][17] ) );
  MUX21X1_RVT U1864 ( .A1(net30566), .A2(net30953), .S0(n158), .Y(n656) );
  IBUFFX4_RVT U1865 ( .A(net30613), .Y(\u_div/PartRem[17][16] ) );
  IBUFFX4_RVT U1866 ( .A(n657), .Y(\u_div/PartRem[17][15] ) );
  MUX21X1_RVT U1867 ( .A1(net30568), .A2(net31003), .S0(n158), .Y(n657) );
  INVX4_RVT U1868 ( .A(n676), .Y(n677) );
  IBUFFX16_RVT U1869 ( .A(\u_div/CryTmp[16][15] ), .Y(n676) );
  INVX1_RVT U1870 ( .A(n658), .Y(\u_div/PartRem[17][14] ) );
  MUX21X1_RVT U1871 ( .A1(net30569), .A2(net31026), .S0(n158), .Y(n658) );
  INVX1_RVT U1872 ( .A(n659), .Y(\u_div/PartRem[17][13] ) );
  MUX21X1_RVT U1873 ( .A1(net30570), .A2(net31048), .S0(net32580), .Y(n659) );
  IBUFFX16_RVT U1874 ( .A(n660), .Y(\u_div/PartRem[17][12] ) );
  MUX21X1_RVT U1875 ( .A1(net30571), .A2(net31070), .S0(net32580), .Y(n660) );
  INVX1_RVT U1876 ( .A(n661), .Y(\u_div/PartRem[17][11] ) );
  MUX21X1_RVT U1877 ( .A1(net30572), .A2(net31090), .S0(net32580), .Y(n661) );
  INVX1_RVT U1878 ( .A(n662), .Y(\u_div/PartRem[17][10] ) );
  MUX21X1_RVT U1879 ( .A1(net30526), .A2(net31109), .S0(net32580), .Y(n662) );
  INVX1_RVT U1880 ( .A(n645), .Y(\u_div/PartRem[17][9] ) );
  MUX21X1_RVT U1881 ( .A1(net30527), .A2(net31127), .S0(net32580), .Y(n645) );
  INVX1_RVT U1882 ( .A(n646), .Y(\u_div/PartRem[17][8] ) );
  INVX1_RVT U1883 ( .A(n647), .Y(\u_div/PartRem[17][7] ) );
  MUX21X1_RVT U1884 ( .A1(net30529), .A2(net31160), .S0(net32580), .Y(n647) );
  INVX1_RVT U1885 ( .A(n648), .Y(\u_div/PartRem[17][6] ) );
  MUX21X1_RVT U1886 ( .A1(net30530), .A2(net31175), .S0(net32580), .Y(n648) );
  INVX1_RVT U1887 ( .A(n650), .Y(\u_div/PartRem[17][4] ) );
  MUX21X1_RVT U1888 ( .A1(net30532), .A2(net31200), .S0(net32580), .Y(n650) );
  MUX21X1_RVT U1889 ( .A1(net30533), .A2(net31211), .S0(n158), .Y(n651) );
  INVX1_RVT U1890 ( .A(n652), .Y(\u_div/PartRem[17][2] ) );
  MUX21X1_RVT U1891 ( .A1(net30562), .A2(net30909), .S0(n158), .Y(n652) );
  MUX21X1_RVT U1892 ( .A1(\u_div/PartRem[16][23] ), .A2(\u_div/SumTmp[15][23] ), .S0(n47), .Y(\u_div/PartRem[15][24] ) );
  INVX1_RVT U1893 ( .A(\u_div/SumTmp[15][22] ), .Y(net30723) );
  INVX0_RVT U1894 ( .A(\u_div/SumTmp[15][21] ), .Y(net30771) );
  INVX0_RVT U1895 ( .A(\u_div/SumTmp[15][20] ), .Y(net30819) );
  INVX0_RVT U1896 ( .A(\u_div/SumTmp[15][19] ), .Y(net30867) );
  INVX0_RVT U1897 ( .A(\u_div/SumTmp[15][18] ), .Y(net30951) );
  IBUFFX16_RVT U1898 ( .A(\u_div/SumTmp[15][16] ), .Y(net31001) );
  INVX0_RVT U1899 ( .A(\u_div/SumTmp[15][15] ), .Y(net31024) );
  INVX0_RVT U1900 ( .A(\u_div/SumTmp[15][14] ), .Y(net31046) );
  INVX0_RVT U1901 ( .A(\u_div/SumTmp[16][13] ), .Y(n665) );
  MUX21X1_RVT U1902 ( .A1(net30662), .A2(net31046), .S0(n51), .Y(net30708) );
  INVX0_RVT U1903 ( .A(\u_div/SumTmp[16][12] ), .Y(n666) );
  INVX0_RVT U1904 ( .A(\u_div/SumTmp[16][11] ), .Y(n667) );
  INVX0_RVT U1905 ( .A(\u_div/SumTmp[16][10] ), .Y(n668) );
  INVX0_RVT U1906 ( .A(\u_div/SumTmp[16][9] ), .Y(n669) );
  INVX0_RVT U1907 ( .A(\u_div/SumTmp[16][8] ), .Y(n670) );
  INVX0_RVT U1908 ( .A(\u_div/SumTmp[16][7] ), .Y(n671) );
  INVX0_RVT U1909 ( .A(\u_div/SumTmp[16][6] ), .Y(n672) );
  INVX0_RVT U1910 ( .A(\u_div/SumTmp[16][5] ), .Y(n673) );
  INVX0_RVT U1911 ( .A(\u_div/SumTmp[16][4] ), .Y(n674) );
  INVX0_RVT U1912 ( .A(\u_div/SumTmp[16][3] ), .Y(n675) );
  INVX0_RVT U1913 ( .A(\u_div/SumTmp[16][2] ), .Y(n664) );
  INVX0_RVT U1914 ( .A(\u_div/SumTmp[16][1] ), .Y(net30917) );
  MUX21X1_RVT U1915 ( .A1(n726), .A2(net31121), .S0(net32542), .Y(net30896) );
  INVX1_RVT U1916 ( .A(net32024), .Y(net32012) );
  INVX1_RVT U1917 ( .A(net30897), .Y(\u_div/PartRem[11][14] ) );
  MUX21X1_RVT U1918 ( .A1(n727), .A2(net31138), .S0(net32544), .Y(net30897) );
  INVX1_RVT U1919 ( .A(b[14]), .Y(net32042) );
  INVX1_RVT U1920 ( .A(net30898), .Y(\u_div/PartRem[11][13] ) );
  MUX21X1_RVT U1921 ( .A1(n728), .A2(net31154), .S0(net32544), .Y(net30898) );
  NBUFFX8_RVT U1922 ( .A(net45939), .Y(net46752) );
  INVX4_RVT U1923 ( .A(n755), .Y(n756) );
  IBUFFX16_RVT U1924 ( .A(\u_div/CryTmp[10][12] ), .Y(n755) );
  INVX4_RVT U1925 ( .A(n750), .Y(n751) );
  INVX1_RVT U1926 ( .A(net30900), .Y(\u_div/PartRem[11][11] ) );
  MUX21X1_RVT U1927 ( .A1(n729), .A2(net31182), .S0(net32542), .Y(net30900) );
  INVX1_RVT U1928 ( .A(net32128), .Y(net32118) );
  INVX1_RVT U1929 ( .A(n744), .Y(n745) );
  INVX1_RVT U1930 ( .A(\u_div/CryTmp[10][11] ), .Y(n744) );
  INVX1_RVT U1931 ( .A(net30901), .Y(\u_div/PartRem[11][10] ) );
  MUX21X1_RVT U1932 ( .A1(n716), .A2(net31194), .S0(net32542), .Y(net30901) );
  INVX1_RVT U1933 ( .A(net32154), .Y(net32144) );
  INVX1_RVT U1934 ( .A(net30855), .Y(\u_div/PartRem[11][9] ) );
  MUX21X1_RVT U1935 ( .A1(n717), .A2(net31205), .S0(net48341), .Y(net30855) );
  INVX1_RVT U1936 ( .A(net30856), .Y(\u_div/PartRem[11][8] ) );
  MUX21X1_RVT U1937 ( .A1(n718), .A2(net30903), .S0(net48341), .Y(net30856) );
  INVX1_RVT U1938 ( .A(net32210), .Y(net32196) );
  INVX1_RVT U1939 ( .A(net30857), .Y(\u_div/PartRem[11][7] ) );
  MUX21X1_RVT U1940 ( .A1(n719), .A2(net30912), .S0(net48341), .Y(net30857) );
  INVX1_RVT U1941 ( .A(net30858), .Y(\u_div/PartRem[11][6] ) );
  MUX21X1_RVT U1942 ( .A1(n720), .A2(net30920), .S0(net48341), .Y(net30858) );
  INVX1_RVT U1943 ( .A(net32264), .Y(net32250) );
  INVX1_RVT U1944 ( .A(net30859), .Y(\u_div/PartRem[11][5] ) );
  MUX21X1_RVT U1945 ( .A1(n721), .A2(net30927), .S0(net48341), .Y(net30859) );
  INVX1_RVT U1946 ( .A(net32300), .Y(net32280) );
  INVX1_RVT U1947 ( .A(net30860), .Y(\u_div/PartRem[11][4] ) );
  MUX21X1_RVT U1948 ( .A1(n722), .A2(net30933), .S0(net48342), .Y(net30860) );
  INVX1_RVT U1949 ( .A(net32324), .Y(net32310) );
  INVX1_RVT U1950 ( .A(net30861), .Y(\u_div/PartRem[11][3] ) );
  MUX21X1_RVT U1951 ( .A1(n723), .A2(net30938), .S0(net48342), .Y(net30861) );
  INVX1_RVT U1952 ( .A(net32352), .Y(net32334) );
  INVX1_RVT U1953 ( .A(net30862), .Y(\u_div/PartRem[11][2] ) );
  MUX21X1_RVT U1954 ( .A1(n724), .A2(net30942), .S0(net48340), .Y(net30862) );
  INVX1_RVT U1955 ( .A(b[2]), .Y(net32362) );
  INVX1_RVT U1956 ( .A(net30891), .Y(\u_div/PartRem[11][1] ) );
  NAND2X0_RVT U1957 ( .A1(net48340), .A2(\*cell*33681/net34095 ), .Y(net30891)
         );
  INVX1_RVT U1958 ( .A(b[0]), .Y(\u_div/CryTmp[11][1] ) );
  INVX0_RVT U1959 ( .A(\u_div/SumTmp[10][15] ), .Y(net31120) );
  INVX0_RVT U1960 ( .A(\u_div/SumTmp[10][14] ), .Y(net31137) );
  INVX0_RVT U1961 ( .A(\u_div/SumTmp[10][13] ), .Y(net31153) );
  INVX0_RVT U1962 ( .A(\u_div/SumTmp[10][12] ), .Y(net31168) );
  MUX21X1_RVT U1963 ( .A1(\u_div/SumTmp[11][11] ), .A2(net45940), .S0(net49094), .Y(net45939) );
  MUX21X1_RVT U1964 ( .A1(net30761), .A2(net31183), .S0(quotient[12]), .Y(n729) );
  INVX1_RVT U1965 ( .A(n716), .Y(\u_div/PartRem[12][9] ) );
  MUX21X1_RVT U1966 ( .A1(net30762), .A2(net31195), .S0(quotient[12]), .Y(n716) );
  INVX1_RVT U1967 ( .A(n717), .Y(\u_div/PartRem[12][8] ) );
  MUX21X1_RVT U1968 ( .A1(net30763), .A2(net31206), .S0(net32548), .Y(n717) );
  INVX1_RVT U1969 ( .A(n718), .Y(\u_div/PartRem[12][7] ) );
  MUX21X1_RVT U1970 ( .A1(net30764), .A2(net30904), .S0(net32548), .Y(n718) );
  INVX1_RVT U1971 ( .A(n719), .Y(\u_div/PartRem[12][6] ) );
  MUX21X1_RVT U1972 ( .A1(net30765), .A2(net30913), .S0(net32548), .Y(n719) );
  INVX1_RVT U1973 ( .A(n720), .Y(\u_div/PartRem[12][5] ) );
  MUX21X1_RVT U1974 ( .A1(net30766), .A2(net30921), .S0(net32548), .Y(n720) );
  INVX1_RVT U1975 ( .A(n721), .Y(\u_div/PartRem[12][4] ) );
  MUX21X1_RVT U1976 ( .A1(net30767), .A2(net30928), .S0(net32548), .Y(n721) );
  INVX1_RVT U1977 ( .A(n722), .Y(\u_div/PartRem[12][3] ) );
  MUX21X1_RVT U1978 ( .A1(net30768), .A2(net30934), .S0(net32548), .Y(n722) );
  INVX1_RVT U1979 ( .A(n723), .Y(\u_div/PartRem[12][2] ) );
  MUX21X1_RVT U1980 ( .A1(net30797), .A2(net30939), .S0(net32548), .Y(n723) );
  INVX1_RVT U1981 ( .A(n724), .Y(\u_div/PartRem[12][1] ) );
  NAND2X0_RVT U1982 ( .A1(net32548), .A2(\*cell*33684/net34105 ), .Y(n724) );
  INVX1_RVT U1983 ( .A(net38336), .Y(net32544) );
  INVX1_RVT U1984 ( .A(net46752), .Y(net30899) );
  AND2X2_RVT U1985 ( .A1(n752), .A2(net46895), .Y(net38336) );
  IBUFFX8_RVT U1986 ( .A(\u_div/PartRem[12][24] ), .Y(n752) );
  MUX21X1_RVT U1987 ( .A1(\u_div/PartRem[13][23] ), .A2(\u_div/SumTmp[12][23] ), .S0(net32548), .Y(\u_div/PartRem[12][24] ) );
  INVX1_RVT U1988 ( .A(\u_div/CryTmp[12][23] ), .Y(n742) );
  IBUFFX4_RVT U1989 ( .A(net30794), .Y(\u_div/PartRem[13][22] ) );
  MUX21X1_RVT U1990 ( .A1(net30748), .A2(net30865), .S0(net42408), .Y(net30794) );
  INVX4_RVT U1991 ( .A(n740), .Y(n741) );
  IBUFFX16_RVT U1992 ( .A(\u_div/CryTmp[12][22] ), .Y(n740) );
  INVX1_RVT U1993 ( .A(net30795), .Y(\u_div/PartRem[13][21] ) );
  INVX1_RVT U1994 ( .A(net30796), .Y(\u_div/PartRem[13][20] ) );
  INVX1_RVT U1995 ( .A(net30798), .Y(\u_div/PartRem[13][19] ) );
  MUX21X1_RVT U1996 ( .A1(n709), .A2(net30999), .S0(net32554), .Y(net30798) );
  INVX4_RVT U1997 ( .A(n759), .Y(n760) );
  IBUFFX16_RVT U1998 ( .A(\u_div/CryTmp[12][19] ), .Y(n759) );
  INVX1_RVT U1999 ( .A(net30799), .Y(\u_div/PartRem[13][18] ) );
  MUX21X1_RVT U2000 ( .A1(n710), .A2(net31022), .S0(net32554), .Y(net30799) );
  IBUFFX4_RVT U2001 ( .A(net30800), .Y(\u_div/PartRem[13][17] ) );
  MUX21X1_RVT U2002 ( .A1(n711), .A2(net31044), .S0(net42408), .Y(net30800) );
  INVX1_RVT U2003 ( .A(net30801), .Y(\u_div/PartRem[13][16] ) );
  MUX21X2_RVT U2004 ( .A1(net30755), .A2(net31066), .S0(net42408), .Y(net30801) );
  INVX1_RVT U2005 ( .A(net30802), .Y(\u_div/PartRem[13][15] ) );
  MUX21X1_RVT U2006 ( .A1(n712), .A2(net31086), .S0(net32554), .Y(net30802) );
  INVX1_RVT U2007 ( .A(net30803), .Y(\u_div/PartRem[13][14] ) );
  MUX21X1_RVT U2008 ( .A1(net30757), .A2(net31105), .S0(net32554), .Y(net30803) );
  INVX1_RVT U2009 ( .A(n715), .Y(\u_div/PartRem[13][13] ) );
  MUX21X1_RVT U2010 ( .A1(net30758), .A2(net31123), .S0(net32554), .Y(n715) );
  MUX21X1_RVT U2011 ( .A1(n696), .A2(net31124), .S0(net47718), .Y(net30758) );
  INVX4_RVT U2012 ( .A(net48671), .Y(net32554) );
  INVX1_RVT U2013 ( .A(net30805), .Y(\u_div/PartRem[13][12] ) );
  MUX21X1_RVT U2014 ( .A1(n713), .A2(net31140), .S0(net32554), .Y(net30805) );
  MUX21X1_RVT U2015 ( .A1(n698), .A2(net31171), .S0(net32554), .Y(net30807) );
  IBUFFX4_RVT U2016 ( .A(net30761), .Y(\u_div/PartRem[13][9] ) );
  MUX21X1_RVT U2017 ( .A1(n699), .A2(n34), .S0(net32554), .Y(net30761) );
  MUX21X1_RVT U2018 ( .A1(n700), .A2(net31196), .S0(net32554), .Y(net30762) );
  INVX1_RVT U2019 ( .A(net30763), .Y(\u_div/PartRem[13][7] ) );
  MUX21X1_RVT U2020 ( .A1(n701), .A2(net31207), .S0(net32554), .Y(net30763) );
  INVX1_RVT U2021 ( .A(net30764), .Y(\u_div/PartRem[13][6] ) );
  MUX21X1_RVT U2022 ( .A1(n702), .A2(net30905), .S0(net32554), .Y(net30764) );
  INVX1_RVT U2023 ( .A(net30765), .Y(\u_div/PartRem[13][5] ) );
  MUX21X1_RVT U2024 ( .A1(n703), .A2(net30914), .S0(net32554), .Y(net30765) );
  INVX1_RVT U2025 ( .A(net30766), .Y(\u_div/PartRem[13][4] ) );
  MUX21X1_RVT U2026 ( .A1(n704), .A2(net30922), .S0(net32554), .Y(net30766) );
  INVX1_RVT U2027 ( .A(net30767), .Y(\u_div/PartRem[13][3] ) );
  MUX21X1_RVT U2028 ( .A1(n705), .A2(net30929), .S0(net32554), .Y(net30767) );
  INVX1_RVT U2029 ( .A(net30768), .Y(\u_div/PartRem[13][2] ) );
  MUX21X1_RVT U2030 ( .A1(n707), .A2(net30935), .S0(net32554), .Y(net30768) );
  INVX1_RVT U2031 ( .A(net30797), .Y(\u_div/PartRem[13][1] ) );
  NAND2X0_RVT U2032 ( .A1(net32554), .A2(\*cell*33687/net34115 ), .Y(net30797)
         );
  INVX4_RVT U2033 ( .A(net38337), .Y(net32548) );
  INVX1_RVT U2034 ( .A(net30841), .Y(\u_div/PartRem[12][22] ) );
  MUX21X1_RVT U2035 ( .A1(net30795), .A2(net30948), .S0(net32548), .Y(net30841) );
  INVX1_RVT U2036 ( .A(net31844), .Y(net31826) );
  INVX1_RVT U2037 ( .A(net30842), .Y(\u_div/PartRem[12][21] ) );
  MUX21X1_RVT U2038 ( .A1(net30796), .A2(net30974), .S0(net32548), .Y(net30842) );
  INVX4_RVT U2039 ( .A(n748), .Y(n749) );
  IBUFFX16_RVT U2040 ( .A(\u_div/CryTmp[11][19] ), .Y(n748) );
  IBUFFX4_RVT U2041 ( .A(net30846), .Y(\u_div/PartRem[12][18] ) );
  MUX21X1_RVT U2042 ( .A1(net30800), .A2(net31043), .S0(quotient[12]), .Y(
        net30846) );
  INVX1_RVT U2043 ( .A(n725), .Y(\u_div/PartRem[12][17] ) );
  MUX21X1_RVT U2044 ( .A1(net30801), .A2(n75), .S0(quotient[12]), .Y(n725) );
  IBUFFX16_RVT U2045 ( .A(\u_div/SumTmp[12][16] ), .Y(net31065) );
  INVX1_RVT U2046 ( .A(net30848), .Y(\u_div/PartRem[12][16] ) );
  MUX21X1_RVT U2047 ( .A1(net30802), .A2(net31085), .S0(quotient[12]), .Y(
        net30848) );
  INVX1_RVT U2048 ( .A(net30849), .Y(\u_div/PartRem[12][15] ) );
  MUX21X1_RVT U2049 ( .A1(net30803), .A2(net31104), .S0(quotient[12]), .Y(
        net30849) );
  MUX21X1_RVT U2050 ( .A1(net45002), .A2(net31122), .S0(n87), .Y(n726) );
  MUX21X1_RVT U2051 ( .A1(net30805), .A2(net31139), .S0(quotient[12]), .Y(n727) );
  INVX4_RVT U2052 ( .A(n753), .Y(n754) );
  IBUFFX16_RVT U2053 ( .A(\u_div/CryTmp[11][12] ), .Y(n753) );
  INVX1_RVT U2054 ( .A(net31922), .Y(net31910) );
  MUX21X1_RVT U2055 ( .A1(\u_div/PartRem[12][23] ), .A2(\u_div/SumTmp[11][23] ), .S0(net32542), .Y(\u_div/PartRem[11][24] ) );
  IBUFFX16_RVT U2056 ( .A(\u_div/SumTmp[11][22] ), .Y(net30947) );
  IBUFFX16_RVT U2057 ( .A(\u_div/SumTmp[12][21] ), .Y(net30948) );
  MUX21X1_RVT U2058 ( .A1(net30841), .A2(net30947), .S0(net32544), .Y(net30946) );
  MUX21X1_RVT U2059 ( .A1(n690), .A2(n731), .S0(net32560), .Y(n706) );
  INVX0_RVT U2060 ( .A(\u_div/SumTmp[13][20] ), .Y(n730) );
  IBUFFX4_RVT U2061 ( .A(n706), .Y(\u_div/PartRem[14][20] ) );
  IBUFFX4_RVT U2062 ( .A(n708), .Y(\u_div/PartRem[14][19] ) );
  MUX21X1_RVT U2063 ( .A1(n691), .A2(n732), .S0(net32560), .Y(n708) );
  IBUFFX4_RVT U2064 ( .A(n709), .Y(\u_div/PartRem[14][18] ) );
  INVX4_RVT U2065 ( .A(n738), .Y(n739) );
  IBUFFX16_RVT U2066 ( .A(\u_div/CryTmp[13][18] ), .Y(n738) );
  INVX1_RVT U2067 ( .A(n710), .Y(\u_div/PartRem[14][17] ) );
  MUX21X1_RVT U2068 ( .A1(n693), .A2(n734), .S0(net32560), .Y(n710) );
  INVX1_RVT U2069 ( .A(n711), .Y(\u_div/PartRem[14][16] ) );
  MUX21X1_RVT U2070 ( .A1(net30708), .A2(n735), .S0(net47718), .Y(n711) );
  INVX1_RVT U2071 ( .A(net30755), .Y(\u_div/PartRem[14][15] ) );
  MUX21X1_RVT U2072 ( .A1(n694), .A2(n736), .S0(net47718), .Y(net30755) );
  INVX1_RVT U2073 ( .A(n712), .Y(\u_div/PartRem[14][14] ) );
  MUX21X1_RVT U2074 ( .A1(n695), .A2(n737), .S0(net47718), .Y(n712) );
  INVX1_RVT U2075 ( .A(net30757), .Y(\u_div/PartRem[14][13] ) );
  INVX1_RVT U2076 ( .A(net30758), .Y(\u_div/PartRem[14][12] ) );
  INVX1_RVT U2077 ( .A(n713), .Y(\u_div/PartRem[14][11] ) );
  MUX21X1_RVT U2078 ( .A1(n697), .A2(net31141), .S0(net47718), .Y(n713) );
  INVX1_RVT U2079 ( .A(n714), .Y(\u_div/PartRem[14][10] ) );
  MUX21X1_RVT U2080 ( .A1(n681), .A2(net31157), .S0(net47718), .Y(n714) );
  INVX1_RVT U2081 ( .A(n698), .Y(\u_div/PartRem[14][9] ) );
  MUX21X1_RVT U2082 ( .A1(n682), .A2(net31172), .S0(net47718), .Y(n698) );
  INVX1_RVT U2083 ( .A(n699), .Y(\u_div/PartRem[14][8] ) );
  MUX21X1_RVT U2084 ( .A1(n683), .A2(net31185), .S0(net47718), .Y(n699) );
  INVX1_RVT U2085 ( .A(n700), .Y(\u_div/PartRem[14][7] ) );
  MUX21X1_RVT U2086 ( .A1(n684), .A2(net31197), .S0(net47718), .Y(n700) );
  MUX21X1_RVT U2087 ( .A1(n685), .A2(net31208), .S0(net32560), .Y(n701) );
  MUX21X1_RVT U2088 ( .A1(n686), .A2(net30906), .S0(net32560), .Y(n702) );
  INVX1_RVT U2089 ( .A(n703), .Y(\u_div/PartRem[14][4] ) );
  MUX21X1_RVT U2090 ( .A1(n687), .A2(net30915), .S0(net32560), .Y(n703) );
  IBUFFX4_RVT U2091 ( .A(n704), .Y(\u_div/PartRem[14][3] ) );
  MUX21X1_RVT U2092 ( .A1(n688), .A2(net30923), .S0(net32560), .Y(n704) );
  IBUFFX4_RVT U2093 ( .A(n705), .Y(\u_div/PartRem[14][2] ) );
  MUX21X1_RVT U2094 ( .A1(n689), .A2(net30930), .S0(net32560), .Y(n705) );
  INVX1_RVT U2095 ( .A(n707), .Y(\u_div/PartRem[14][1] ) );
  NAND2X0_RVT U2096 ( .A1(net32560), .A2(\*cell*33690/net34125 ), .Y(n707) );
  INVX1_RVT U2097 ( .A(net48671), .Y(net42408) );
  MUX21X1_RVT U2098 ( .A1(net30658), .A2(net30951), .S0(n48), .Y(n690) );
  INVX0_RVT U2099 ( .A(\u_div/SumTmp[14][19] ), .Y(n731) );
  INVX1_RVT U2100 ( .A(n690), .Y(\u_div/PartRem[15][19] ) );
  IBUFFX16_RVT U2101 ( .A(n691), .Y(\u_div/PartRem[15][18] ) );
  MUX21X1_RVT U2102 ( .A1(net30660), .A2(net31001), .S0(n59), .Y(n692) );
  MUX21X1_RVT U2103 ( .A1(net30661), .A2(net31024), .S0(n55), .Y(n693) );
  INVX1_RVT U2104 ( .A(net30708), .Y(\u_div/PartRem[15][15] ) );
  INVX1_RVT U2105 ( .A(n694), .Y(\u_div/PartRem[15][14] ) );
  MUX21X1_RVT U2106 ( .A1(net30663), .A2(net31068), .S0(n48), .Y(n694) );
  INVX1_RVT U2107 ( .A(n695), .Y(\u_div/PartRem[15][13] ) );
  MUX21X2_RVT U2108 ( .A1(net30664), .A2(net31088), .S0(n46), .Y(n695) );
  INVX2_RVT U2109 ( .A(net42405), .Y(net42406) );
  IBUFFX16_RVT U2110 ( .A(\u_div/CryTmp[14][12] ), .Y(net42405) );
  INVX1_RVT U2111 ( .A(n696), .Y(\u_div/PartRem[15][11] ) );
  MUX21X1_RVT U2112 ( .A1(net30666), .A2(net31125), .S0(n52), .Y(n696) );
  INVX1_RVT U2113 ( .A(n697), .Y(\u_div/PartRem[15][10] ) );
  MUX21X1_RVT U2114 ( .A1(net30620), .A2(net31142), .S0(n50), .Y(n697) );
  INVX1_RVT U2115 ( .A(n681), .Y(\u_div/PartRem[15][9] ) );
  MUX21X1_RVT U2116 ( .A1(net30621), .A2(net31158), .S0(n49), .Y(n681) );
  INVX1_RVT U2117 ( .A(n682), .Y(\u_div/PartRem[15][8] ) );
  MUX21X1_RVT U2118 ( .A1(net30622), .A2(net31173), .S0(n45), .Y(n682) );
  INVX1_RVT U2119 ( .A(n683), .Y(\u_div/PartRem[15][7] ) );
  MUX21X1_RVT U2120 ( .A1(net30623), .A2(net31186), .S0(n57), .Y(n683) );
  INVX1_RVT U2121 ( .A(n684), .Y(\u_div/PartRem[15][6] ) );
  MUX21X1_RVT U2122 ( .A1(net30624), .A2(net31198), .S0(n54), .Y(n684) );
  INVX1_RVT U2123 ( .A(n685), .Y(\u_div/PartRem[15][5] ) );
  MUX21X1_RVT U2124 ( .A1(net30625), .A2(net31209), .S0(n51), .Y(n685) );
  INVX1_RVT U2125 ( .A(n686), .Y(\u_div/PartRem[15][4] ) );
  MUX21X2_RVT U2126 ( .A1(net30626), .A2(net30907), .S0(n49), .Y(n686) );
  INVX1_RVT U2127 ( .A(n687), .Y(\u_div/PartRem[15][3] ) );
  INVX1_RVT U2128 ( .A(n688), .Y(\u_div/PartRem[15][2] ) );
  MUX21X1_RVT U2129 ( .A1(net30656), .A2(net30924), .S0(n46), .Y(n688) );
  INVX4_RVT U2130 ( .A(n757), .Y(n758) );
  IBUFFX4_RVT U2131 ( .A(\u_div/PartRem[15][1] ), .Y(n757) );
  INVX0_RVT U2132 ( .A(n689), .Y(\u_div/PartRem[15][1] ) );
  NAND2X0_RVT U2133 ( .A1(n59), .A2(\*cell*33693/net34135 ), .Y(n689) );
  INVX0_RVT U2134 ( .A(\u_div/SumTmp[14][18] ), .Y(n732) );
  INVX0_RVT U2135 ( .A(\u_div/SumTmp[14][17] ), .Y(n733) );
  INVX0_RVT U2136 ( .A(\u_div/SumTmp[14][16] ), .Y(n734) );
  INVX0_RVT U2137 ( .A(\u_div/SumTmp[14][15] ), .Y(n735) );
  INVX0_RVT U2138 ( .A(\u_div/SumTmp[14][14] ), .Y(n736) );
  IBUFFX4_RVT U2139 ( .A(\u_div/SumTmp[14][13] ), .Y(n737) );
  INVX0_RVT U2140 ( .A(\u_div/SumTmp[14][12] ), .Y(net31106) );
  MUX21X1_RVT U2141 ( .A1(net29739), .A2(net29740), .S0(net32530), .Y(n761) );
  INVX0_RVT U2142 ( .A(\u_div/SumTmp[8][19] ), .Y(net29738) );
  IBUFFX4_RVT U2143 ( .A(n761), .Y(\u_div/PartRem[9][19] ) );
  IBUFFX4_RVT U2144 ( .A(net29611), .Y(\u_div/PartRem[9][18] ) );
  MUX21X1_RVT U2145 ( .A1(net29797), .A2(net29798), .S0(net32530), .Y(net29611) );
  IBUFFX4_RVT U2146 ( .A(net29612), .Y(\u_div/PartRem[9][17] ) );
  MUX21X1_RVT U2147 ( .A1(net29945), .A2(net29946), .S0(net32530), .Y(net29612) );
  IBUFFX4_RVT U2148 ( .A(net29613), .Y(\u_div/PartRem[9][16] ) );
  MUX21X1_RVT U2149 ( .A1(net30337), .A2(net30338), .S0(net32530), .Y(net29613) );
  IBUFFX4_RVT U2150 ( .A(net29614), .Y(\u_div/PartRem[9][15] ) );
  MUX21X1_RVT U2151 ( .A1(net30347), .A2(net30348), .S0(net32530), .Y(net29614) );
  IBUFFX4_RVT U2152 ( .A(net49255), .Y(\u_div/PartRem[9][14] ) );
  INVX4_RVT U2153 ( .A(net49254), .Y(net49255) );
  INVX4_RVT U2154 ( .A(n769), .Y(n770) );
  IBUFFX16_RVT U2155 ( .A(\u_div/CryTmp[8][14] ), .Y(n769) );
  INVX1_RVT U2156 ( .A(net29616), .Y(\u_div/PartRem[9][13] ) );
  MUX21X1_RVT U2157 ( .A1(net30367), .A2(net30368), .S0(net32530), .Y(net29616) );
  INVX1_RVT U2158 ( .A(net32076), .Y(net32068) );
  INVX1_RVT U2159 ( .A(net29617), .Y(\u_div/PartRem[9][12] ) );
  MUX21X1_RVT U2160 ( .A1(net30377), .A2(net30378), .S0(net46550), .Y(net29617) );
  INVX1_RVT U2161 ( .A(net29618), .Y(\u_div/PartRem[9][11] ) );
  MUX21X1_RVT U2162 ( .A1(net30387), .A2(net30388), .S0(net46550), .Y(net29618) );
  IBUFFX16_RVT U2163 ( .A(n773), .Y(n774) );
  INVX2_RVT U2164 ( .A(net29619), .Y(\u_div/PartRem[9][10] ) );
  INVX1_RVT U2165 ( .A(net29598), .Y(\u_div/PartRem[9][9] ) );
  MUX21X1_RVT U2166 ( .A1(net30407), .A2(net30408), .S0(net46550), .Y(net29598) );
  INVX1_RVT U2167 ( .A(net29599), .Y(\u_div/PartRem[9][8] ) );
  MUX21X1_RVT U2168 ( .A1(net30417), .A2(net30418), .S0(net46550), .Y(net29599) );
  INVX1_RVT U2169 ( .A(net29600), .Y(\u_div/PartRem[9][7] ) );
  MUX21X1_RVT U2170 ( .A1(net30427), .A2(net30428), .S0(net46550), .Y(net29600) );
  MUX21X1_RVT U2171 ( .A1(net30447), .A2(net30448), .S0(net46550), .Y(net29602) );
  MUX21X1_RVT U2172 ( .A1(net30457), .A2(net30458), .S0(net46550), .Y(net29603) );
  INVX1_RVT U2173 ( .A(net29605), .Y(\u_div/PartRem[9][2] ) );
  MUX21X1_RVT U2174 ( .A1(net30477), .A2(net30478), .S0(net32530), .Y(net29605) );
  INVX1_RVT U2175 ( .A(net29609), .Y(\u_div/PartRem[9][1] ) );
  NAND2X0_RVT U2176 ( .A1(net32530), .A2(\*cell*33726/net34245 ), .Y(net29609)
         );
  MUX21X1_RVT U2177 ( .A1(net30467), .A2(net30468), .S0(net46550), .Y(net29604) );
  MUX21X1_RVT U2178 ( .A1(net29633), .A2(net29737), .S0(net46859), .Y(net29658) );
  MUX21X1_RVT U2179 ( .A1(n764), .A2(n765), .S0(net32538), .Y(net29739) );
  INVX0_RVT U2180 ( .A(\u_div/SumTmp[9][18] ), .Y(net29740) );
  INVX1_RVT U2181 ( .A(net29739), .Y(\u_div/PartRem[10][18] ) );
  INVX1_RVT U2182 ( .A(net29797), .Y(\u_div/PartRem[10][17] ) );
  MUX21X1_RVT U2183 ( .A1(net30895), .A2(net31102), .S0(net32538), .Y(net29797) );
  INVX1_RVT U2184 ( .A(net29945), .Y(\u_div/PartRem[10][16] ) );
  MUX21X1_RVT U2185 ( .A1(net30896), .A2(net31120), .S0(net32538), .Y(net29945) );
  INVX1_RVT U2186 ( .A(net30337), .Y(\u_div/PartRem[10][15] ) );
  MUX21X1_RVT U2187 ( .A1(net30897), .A2(net31137), .S0(net32538), .Y(net30337) );
  INVX1_RVT U2188 ( .A(net30347), .Y(\u_div/PartRem[10][14] ) );
  MUX21X1_RVT U2189 ( .A1(net30898), .A2(net31153), .S0(net32538), .Y(net30347) );
  INVX1_RVT U2190 ( .A(net30357), .Y(\u_div/PartRem[10][13] ) );
  MUX21X1_RVT U2191 ( .A1(net30899), .A2(net31168), .S0(net32538), .Y(net30357) );
  INVX1_RVT U2192 ( .A(net30367), .Y(\u_div/PartRem[10][12] ) );
  MUX21X1_RVT U2193 ( .A1(net30900), .A2(net31181), .S0(net32538), .Y(net30367) );
  INVX1_RVT U2194 ( .A(net30377), .Y(\u_div/PartRem[10][11] ) );
  MUX21X1_RVT U2195 ( .A1(net30901), .A2(net31193), .S0(net32538), .Y(net30377) );
  INVX1_RVT U2196 ( .A(net30387), .Y(\u_div/PartRem[10][10] ) );
  MUX21X1_RVT U2197 ( .A1(net30855), .A2(net31204), .S0(net32536), .Y(net30387) );
  INVX1_RVT U2198 ( .A(net30397), .Y(\u_div/PartRem[10][9] ) );
  MUX21X1_RVT U2199 ( .A1(net30856), .A2(net30902), .S0(net32536), .Y(net30397) );
  MUX21X1_RVT U2200 ( .A1(net30857), .A2(net30911), .S0(net32536), .Y(net30407) );
  MUX21X1_RVT U2201 ( .A1(net30858), .A2(net30919), .S0(net32536), .Y(net30417) );
  INVX1_RVT U2202 ( .A(net30427), .Y(\u_div/PartRem[10][6] ) );
  MUX21X1_RVT U2203 ( .A1(net30859), .A2(net30926), .S0(net32536), .Y(net30427) );
  INVX1_RVT U2204 ( .A(n762), .Y(\u_div/PartRem[10][5] ) );
  MUX21X1_RVT U2205 ( .A1(net30860), .A2(net30932), .S0(net32536), .Y(n762) );
  IBUFFX16_RVT U2206 ( .A(\u_div/CryTmp[9][5] ), .Y(n767) );
  INVX1_RVT U2207 ( .A(net30447), .Y(\u_div/PartRem[10][4] ) );
  MUX21X1_RVT U2208 ( .A1(net30861), .A2(net30937), .S0(net32536), .Y(net30447) );
  INVX1_RVT U2209 ( .A(net30457), .Y(\u_div/PartRem[10][3] ) );
  MUX21X1_RVT U2210 ( .A1(net30862), .A2(net30941), .S0(net32536), .Y(net30457) );
  IBUFFX2_RVT U2211 ( .A(net30467), .Y(\u_div/PartRem[10][2] ) );
  INVX1_RVT U2212 ( .A(net30477), .Y(\u_div/PartRem[10][1] ) );
  NAND2X0_RVT U2213 ( .A1(net32538), .A2(\*cell*33690/net34125 ), .Y(net30477)
         );
  INVX4_RVT U2214 ( .A(net45541), .Y(net32530) );
  INVX0_RVT U2215 ( .A(\u_div/SumTmp[9][17] ), .Y(net29798) );
  INVX0_RVT U2216 ( .A(\u_div/SumTmp[9][16] ), .Y(net29946) );
  INVX0_RVT U2217 ( .A(\u_div/SumTmp[9][15] ), .Y(net30338) );
  INVX0_RVT U2218 ( .A(\u_div/SumTmp[9][14] ), .Y(net30348) );
  IBUFFX16_RVT U2219 ( .A(\u_div/SumTmp[9][13] ), .Y(net30358) );
  INVX0_RVT U2220 ( .A(\u_div/SumTmp[9][12] ), .Y(net30368) );
  INVX0_RVT U2221 ( .A(\u_div/SumTmp[9][11] ), .Y(net30378) );
  INVX0_RVT U2222 ( .A(\u_div/SumTmp[9][10] ), .Y(net30388) );
  INVX0_RVT U2223 ( .A(\u_div/SumTmp[9][9] ), .Y(net30398) );
  INVX0_RVT U2224 ( .A(\u_div/SumTmp[9][8] ), .Y(net30408) );
  INVX0_RVT U2225 ( .A(\u_div/SumTmp[9][7] ), .Y(net30418) );
  INVX0_RVT U2226 ( .A(\u_div/SumTmp[9][6] ), .Y(net30428) );
  INVX0_RVT U2227 ( .A(\u_div/SumTmp[9][5] ), .Y(n763) );
  INVX0_RVT U2228 ( .A(\u_div/SumTmp[10][4] ), .Y(net30932) );
  INVX0_RVT U2229 ( .A(n766), .Y(net32536) );
  MUX21X1_RVT U2230 ( .A1(n762), .A2(n763), .S0(net46550), .Y(net29601) );
  NOR2X1_RVT U2231 ( .A1(\u_div/PartRem[11][24] ), .A2(\u_div/CryTmp[10][24] ), 
        .Y(n766) );
  INVX1_RVT U2232 ( .A(net30946), .Y(\u_div/PartRem[11][23] ) );
  INVX1_RVT U2233 ( .A(net30888), .Y(\u_div/PartRem[11][22] ) );
  INVX1_RVT U2234 ( .A(net30889), .Y(\u_div/PartRem[11][21] ) );
  INVX1_RVT U2235 ( .A(net30892), .Y(\u_div/PartRem[11][19] ) );
  INVX1_RVT U2236 ( .A(net30893), .Y(\u_div/PartRem[11][18] ) );
  INVX1_RVT U2237 ( .A(n764), .Y(\u_div/PartRem[11][17] ) );
  MUX21X1_RVT U2238 ( .A1(net30848), .A2(net31084), .S0(net32544), .Y(n764) );
  MUX21X1_RVT U2239 ( .A1(net30849), .A2(net31103), .S0(net32542), .Y(net30895) );
  INVX4_RVT U2240 ( .A(n766), .Y(net32538) );
  MUX21X1_RVT U2241 ( .A1(\u_div/PartRem[11][23] ), .A2(\u_div/SumTmp[10][23] ), .S0(net32536), .Y(\u_div/PartRem[10][24] ) );
  INVX1_RVT U2242 ( .A(\u_div/SumTmp[10][22] ), .Y(net30972) );
  INVX0_RVT U2243 ( .A(\u_div/SumTmp[10][21] ), .Y(net30996) );
  INVX0_RVT U2244 ( .A(\u_div/SumTmp[10][20] ), .Y(net31019) );
  INVX0_RVT U2245 ( .A(\u_div/SumTmp[10][19] ), .Y(net31041) );
  INVX0_RVT U2246 ( .A(\u_div/SumTmp[10][18] ), .Y(net31063) );
  INVX0_RVT U2247 ( .A(\u_div/SumTmp[10][17] ), .Y(n765) );
  INVX0_RVT U2248 ( .A(\u_div/SumTmp[10][16] ), .Y(net31102) );
  INVX0_RVT U2249 ( .A(net42548), .Y(net45600) );
  INVX1_RVT U2250 ( .A(n842), .Y(net42548) );
  MUX21X1_RVT U2251 ( .A1(n822), .A2(net30351), .S0(net45604), .Y(net29801) );
  MUX21X1_RVT U2252 ( .A1(n809), .A2(net29940), .S0(net50726), .Y(net29741) );
  INVX1_RVT U2253 ( .A(net29742), .Y(\u_div/PartRem[4][21] ) );
  MUX21X1_RVT U2254 ( .A1(n810), .A2(net30332), .S0(net50726), .Y(net29742) );
  INVX1_RVT U2255 ( .A(net29743), .Y(\u_div/PartRem[4][20] ) );
  MUX21X1_RVT U2256 ( .A1(n812), .A2(net30342), .S0(net50726), .Y(net29743) );
  MUX21X1_RVT U2257 ( .A1(n813), .A2(net30352), .S0(net42034), .Y(n822) );
  INVX1_RVT U2258 ( .A(net29746), .Y(\u_div/PartRem[4][18] ) );
  MUX21X1_RVT U2259 ( .A1(n814), .A2(net30362), .S0(net42034), .Y(net29746) );
  INVX1_RVT U2260 ( .A(net29747), .Y(\u_div/PartRem[4][17] ) );
  MUX21X1_RVT U2261 ( .A1(n815), .A2(net30372), .S0(net42034), .Y(net29747) );
  INVX1_RVT U2262 ( .A(net31972), .Y(net31964) );
  INVX1_RVT U2263 ( .A(net29748), .Y(\u_div/PartRem[4][16] ) );
  MUX21X1_RVT U2264 ( .A1(n816), .A2(net30382), .S0(net42034), .Y(net29748) );
  INVX1_RVT U2265 ( .A(net31998), .Y(net31986) );
  INVX1_RVT U2266 ( .A(net29749), .Y(\u_div/PartRem[4][15] ) );
  MUX21X1_RVT U2267 ( .A1(n817), .A2(net30392), .S0(net42034), .Y(net29749) );
  INVX1_RVT U2268 ( .A(net29750), .Y(\u_div/PartRem[4][14] ) );
  MUX21X1_RVT U2269 ( .A1(n818), .A2(net30402), .S0(net42034), .Y(net29750) );
  MUX21X1_RVT U2270 ( .A1(n819), .A2(net30412), .S0(net40598), .Y(net29751) );
  MUX21X1_RVT U2271 ( .A1(n820), .A2(net30422), .S0(net42034), .Y(net29752) );
  INVX1_RVT U2272 ( .A(net29753), .Y(\u_div/PartRem[4][11] ) );
  MUX21X1_RVT U2273 ( .A1(n821), .A2(net30432), .S0(net50726), .Y(net29753) );
  INVX1_RVT U2274 ( .A(n823), .Y(\u_div/PartRem[4][10] ) );
  MUX21X1_RVT U2275 ( .A1(net29698), .A2(net46608), .S0(net50726), .Y(n823) );
  MUX21X1_RVT U2276 ( .A1(net29672), .A2(net30443), .S0(net49625), .Y(net29698) );
  INVX1_RVT U2277 ( .A(net29726), .Y(\u_div/PartRem[4][9] ) );
  MUX21X1_RVT U2278 ( .A1(n803), .A2(net45229), .S0(net50726), .Y(net29726) );
  INVX1_RVT U2279 ( .A(net29727), .Y(\u_div/PartRem[4][8] ) );
  INVX1_RVT U2280 ( .A(net29728), .Y(\u_div/PartRem[4][7] ) );
  MUX21X1_RVT U2281 ( .A1(n805), .A2(net30472), .S0(net42034), .Y(net29728) );
  INVX1_RVT U2282 ( .A(n843), .Y(n844) );
  INVX1_RVT U2283 ( .A(net29730), .Y(\u_div/PartRem[4][5] ) );
  MUX21X1_RVT U2284 ( .A1(n806), .A2(net30297), .S0(net50726), .Y(net29730) );
  INVX1_RVT U2285 ( .A(net29731), .Y(\u_div/PartRem[4][4] ) );
  MUX21X1_RVT U2286 ( .A1(n807), .A2(net30305), .S0(net50726), .Y(net29731) );
  INVX1_RVT U2287 ( .A(net29732), .Y(\u_div/PartRem[4][3] ) );
  MUX21X1_RVT U2288 ( .A1(n808), .A2(net30312), .S0(net50726), .Y(net29732) );
  INVX1_RVT U2289 ( .A(net29733), .Y(\u_div/PartRem[4][2] ) );
  MUX21X1_RVT U2290 ( .A1(n811), .A2(net30318), .S0(net50726), .Y(net29733) );
  INVX1_RVT U2291 ( .A(net29744), .Y(\u_div/PartRem[4][1] ) );
  NAND2X0_RVT U2292 ( .A1(net50726), .A2(\u_div/SumTmp[5][0] ), .Y(net29744)
         );
  INVX1_RVT U2293 ( .A(n810), .Y(\u_div/PartRem[5][20] ) );
  MUX21X1_RVT U2294 ( .A1(n793), .A2(n825), .S0(net49601), .Y(n810) );
  MUX21X1_RVT U2295 ( .A1(n794), .A2(n826), .S0(net49611), .Y(n812) );
  INVX1_RVT U2296 ( .A(n813), .Y(\u_div/PartRem[5][18] ) );
  MUX21X1_RVT U2297 ( .A1(n795), .A2(n827), .S0(net44755), .Y(n813) );
  INVX1_RVT U2298 ( .A(n814), .Y(\u_div/PartRem[5][17] ) );
  MUX21X1_RVT U2299 ( .A1(n796), .A2(n828), .S0(net44755), .Y(n814) );
  INVX1_RVT U2300 ( .A(n815), .Y(\u_div/PartRem[5][16] ) );
  MUX21X1_RVT U2301 ( .A1(n797), .A2(n829), .S0(quotient[5]), .Y(n815) );
  INVX1_RVT U2302 ( .A(n816), .Y(\u_div/PartRem[5][15] ) );
  INVX1_RVT U2303 ( .A(n817), .Y(\u_div/PartRem[5][14] ) );
  MUX21X1_RVT U2304 ( .A1(n799), .A2(n831), .S0(net44755), .Y(n817) );
  INVX1_RVT U2305 ( .A(n818), .Y(\u_div/PartRem[5][13] ) );
  MUX21X1_RVT U2306 ( .A1(n800), .A2(n832), .S0(net44755), .Y(n818) );
  INVX1_RVT U2307 ( .A(n819), .Y(\u_div/PartRem[5][12] ) );
  MUX21X1_RVT U2308 ( .A1(n801), .A2(n833), .S0(net44755), .Y(n819) );
  INVX1_RVT U2309 ( .A(n820), .Y(\u_div/PartRem[5][11] ) );
  MUX21X1_RVT U2310 ( .A1(n802), .A2(n834), .S0(n128), .Y(n820) );
  INVX1_RVT U2311 ( .A(n821), .Y(\u_div/PartRem[5][10] ) );
  MUX21X1_RVT U2312 ( .A1(net29671), .A2(net30433), .S0(net32506), .Y(n821) );
  INVX1_RVT U2313 ( .A(net29698), .Y(\u_div/PartRem[5][9] ) );
  INVX1_RVT U2314 ( .A(n803), .Y(\u_div/PartRem[5][8] ) );
  MUX21X1_RVT U2315 ( .A1(n787), .A2(net30453), .S0(net49611), .Y(n803) );
  INVX1_RVT U2316 ( .A(n805), .Y(\u_div/PartRem[5][6] ) );
  MUX21X1_RVT U2317 ( .A1(n788), .A2(net30473), .S0(net44755), .Y(n805) );
  MUX21X1_RVT U2318 ( .A1(n784), .A2(net30289), .S0(net45257), .Y(net29676) );
  INVX1_RVT U2319 ( .A(n806), .Y(\u_div/PartRem[5][4] ) );
  MUX21X1_RVT U2320 ( .A1(n789), .A2(net30298), .S0(quotient[5]), .Y(n806) );
  INVX1_RVT U2321 ( .A(n807), .Y(\u_div/PartRem[5][3] ) );
  MUX21X1_RVT U2322 ( .A1(n790), .A2(net30306), .S0(quotient[5]), .Y(n807) );
  INVX1_RVT U2323 ( .A(n808), .Y(\u_div/PartRem[5][2] ) );
  MUX21X1_RVT U2324 ( .A1(n792), .A2(net30313), .S0(net44755), .Y(n808) );
  INVX1_RVT U2325 ( .A(n811), .Y(\u_div/PartRem[5][1] ) );
  NAND2X0_RVT U2326 ( .A1(net44755), .A2(\u_div/SumTmp[5][0] ), .Y(n811) );
  MUX21X1_RVT U2327 ( .A1(n873), .A2(\u_div/SumTmp[4][22] ), .S0(n176), .Y(
        net38274) );
  INVX2_RVT U2328 ( .A(net29685), .Y(\u_div/PartRem[6][21] ) );
  INVX1_RVT U2329 ( .A(n791), .Y(\u_div/PartRem[6][20] ) );
  MUX21X1_RVT U2330 ( .A1(net29661), .A2(net29942), .S0(net45257), .Y(n791) );
  MUX21X1_RVT U2331 ( .A1(net29662), .A2(net30334), .S0(net45257), .Y(n793) );
  INVX1_RVT U2332 ( .A(n794), .Y(\u_div/PartRem[6][18] ) );
  MUX21X1_RVT U2333 ( .A1(net29663), .A2(net30344), .S0(net45257), .Y(n794) );
  INVX1_RVT U2334 ( .A(n795), .Y(\u_div/PartRem[6][17] ) );
  INVX1_RVT U2335 ( .A(n796), .Y(\u_div/PartRem[6][16] ) );
  MUX21X1_RVT U2336 ( .A1(net29665), .A2(net30364), .S0(net45257), .Y(n796) );
  INVX1_RVT U2337 ( .A(n798), .Y(\u_div/PartRem[6][14] ) );
  INVX1_RVT U2338 ( .A(n799), .Y(\u_div/PartRem[6][13] ) );
  INVX1_RVT U2339 ( .A(n800), .Y(\u_div/PartRem[6][12] ) );
  MUX21X1_RVT U2340 ( .A1(net29669), .A2(net30404), .S0(net45257), .Y(n800) );
  INVX1_RVT U2341 ( .A(n801), .Y(\u_div/PartRem[6][11] ) );
  MUX21X1_RVT U2342 ( .A1(net29670), .A2(net30414), .S0(net45257), .Y(n801) );
  MUX21X1_RVT U2343 ( .A1(\u_div/SumTmp[6][8] ), .A2(\u_div/PartRem[7][8] ), 
        .S0(net52013), .Y(net52003) );
  MUX21X1_RVT U2344 ( .A1(\u_div/SumTmp[6][7] ), .A2(\u_div/PartRem[7][7] ), 
        .S0(net45737), .Y(net52000) );
  INVX1_RVT U2345 ( .A(n788), .Y(\u_div/PartRem[6][5] ) );
  MUX21X1_RVT U2346 ( .A1(n783), .A2(net30474), .S0(net45257), .Y(n788) );
  INVX1_RVT U2347 ( .A(net29676), .Y(\u_div/PartRem[6][4] ) );
  INVX1_RVT U2348 ( .A(n789), .Y(\u_div/PartRem[6][3] ) );
  MUX21X2_RVT U2349 ( .A1(n785), .A2(net30299), .S0(net40656), .Y(n789) );
  INVX1_RVT U2350 ( .A(n790), .Y(\u_div/PartRem[6][2] ) );
  MUX21X1_RVT U2351 ( .A1(n786), .A2(net30307), .S0(net45257), .Y(n790) );
  INVX1_RVT U2352 ( .A(n792), .Y(\u_div/PartRem[6][1] ) );
  NAND2X0_RVT U2353 ( .A1(net45257), .A2(\*cell*33717/net34215 ), .Y(n792) );
  INVX0_RVT U2354 ( .A(n787), .Y(n874) );
  INVX0_RVT U2355 ( .A(\u_div/SumTmp[5][19] ), .Y(n825) );
  INVX0_RVT U2356 ( .A(\u_div/SumTmp[5][18] ), .Y(n826) );
  INVX0_RVT U2357 ( .A(\u_div/SumTmp[5][17] ), .Y(n827) );
  INVX0_RVT U2358 ( .A(\u_div/SumTmp[5][16] ), .Y(n828) );
  INVX0_RVT U2359 ( .A(\u_div/SumTmp[5][15] ), .Y(n829) );
  INVX0_RVT U2360 ( .A(\u_div/SumTmp[5][13] ), .Y(n831) );
  INVX0_RVT U2361 ( .A(\u_div/SumTmp[5][12] ), .Y(n832) );
  INVX0_RVT U2362 ( .A(\u_div/SumTmp[5][11] ), .Y(n833) );
  INVX0_RVT U2363 ( .A(\u_div/SumTmp[5][10] ), .Y(n834) );
  INVX1_RVT U2364 ( .A(n782), .Y(\u_div/PartRem[7][9] ) );
  MUX21X1_RVT U2365 ( .A1(n777), .A2(n835), .S0(net46768), .Y(n782) );
  INVX2_RVT U2366 ( .A(net29646), .Y(\u_div/PartRem[7][8] ) );
  INVX2_RVT U2367 ( .A(net29647), .Y(\u_div/PartRem[7][7] ) );
  INVX1_RVT U2368 ( .A(net29649), .Y(\u_div/PartRem[7][5] ) );
  MUX21X1_RVT U2369 ( .A1(n778), .A2(net30465), .S0(net46768), .Y(net29649) );
  INVX1_RVT U2370 ( .A(n783), .Y(\u_div/PartRem[7][4] ) );
  MUX21X1_RVT U2371 ( .A1(n779), .A2(net30475), .S0(net46768), .Y(n783) );
  INVX1_RVT U2372 ( .A(n785), .Y(\u_div/PartRem[7][2] ) );
  MUX21X1_RVT U2373 ( .A1(n781), .A2(net30300), .S0(net46859), .Y(n785) );
  INVX1_RVT U2374 ( .A(n786), .Y(\u_div/PartRem[7][1] ) );
  NAND2X0_RVT U2375 ( .A1(net46768), .A2(\*cell*33720/net34225 ), .Y(n786) );
  INVX2_RVT U2376 ( .A(net29648), .Y(\u_div/PartRem[7][6] ) );
  MUX21X1_RVT U2377 ( .A1(net29600), .A2(net30426), .S0(net40719), .Y(n777) );
  INVX0_RVT U2378 ( .A(\u_div/SumTmp[7][8] ), .Y(n835) );
  INVX1_RVT U2379 ( .A(n777), .Y(\u_div/PartRem[8][8] ) );
  MUX21X1_RVT U2380 ( .A1(\u_div/SumTmp[8][6] ), .A2(\u_div/PartRem[9][6] ), 
        .S0(net40717), .Y(net40783) );
  INVX1_RVT U2381 ( .A(net29623), .Y(\u_div/PartRem[8][6] ) );
  MUX21X1_RVT U2382 ( .A1(net29602), .A2(net30446), .S0(net40719), .Y(net29623) );
  INVX1_RVT U2383 ( .A(net29624), .Y(\u_div/PartRem[8][5] ) );
  MUX21X1_RVT U2384 ( .A1(net29603), .A2(net30456), .S0(net40719), .Y(net29624) );
  INVX1_RVT U2385 ( .A(n778), .Y(\u_div/PartRem[8][4] ) );
  MUX21X1_RVT U2386 ( .A1(net29604), .A2(net30466), .S0(net40719), .Y(n778) );
  INVX1_RVT U2387 ( .A(n779), .Y(\u_div/PartRem[8][3] ) );
  MUX21X1_RVT U2388 ( .A1(net29605), .A2(net30476), .S0(net40719), .Y(n779) );
  NAND2X0_RVT U2389 ( .A1(net40724), .A2(\*cell*33723/net34235 ), .Y(n781) );
  INVX1_RVT U2390 ( .A(net38347), .Y(net46768) );
  NOR2X1_RVT U2391 ( .A1(\u_div/PartRem[8][24] ), .A2(\u_div/CryTmp[7][24] ), 
        .Y(net38347) );
  MUX21X1_RVT U2392 ( .A1(\u_div/PartRem[9][23] ), .A2(\u_div/SumTmp[8][23] ), 
        .S0(net40720), .Y(\u_div/PartRem[8][24] ) );
  IBUFFX4_RVT U2393 ( .A(net29628), .Y(\u_div/PartRem[9][23] ) );
  INVX1_RVT U2394 ( .A(net29606), .Y(\u_div/PartRem[9][22] ) );
  MUX21X1_RVT U2395 ( .A1(net29655), .A2(net51612), .S0(net32530), .Y(net29606) );
  MUX21X1_RVT U2396 ( .A1(net29682), .A2(net29683), .S0(net32530), .Y(n775) );
  IBUFFX4_RVT U2397 ( .A(n776), .Y(\u_div/PartRem[9][20] ) );
  MUX21X1_RVT U2398 ( .A1(net29710), .A2(net29711), .S0(net32530), .Y(n776) );
  INVX1_RVT U2399 ( .A(net29653), .Y(\u_div/PartRem[8][23] ) );
  INVX1_RVT U2400 ( .A(net29631), .Y(\u_div/PartRem[8][22] ) );
  MUX21X1_RVT U2401 ( .A1(n775), .A2(net29681), .S0(net40720), .Y(net29631) );
  INVX4_RVT U2402 ( .A(net29632), .Y(n855) );
  MUX21X2_RVT U2403 ( .A1(n776), .A2(net29709), .S0(net40718), .Y(net29632) );
  INVX16_RVT U2404 ( .A(net29635), .Y(\u_div/PartRem[8][19] ) );
  MUX21X2_RVT U2405 ( .A1(net29611), .A2(net29796), .S0(net40718), .Y(net29635) );
  NAND3X0_RVT U2406 ( .A1(n839), .A2(n838), .A3(n837), .Y(
        \u_div/CryTmp[7][19] ) );
  NAND2X0_RVT U2407 ( .A1(net31940), .A2(\u_div/PartRem[8][18] ), .Y(n839) );
  INVX2_RVT U2408 ( .A(n260), .Y(\u_div/PartRem[8][18] ) );
  NAND2X0_RVT U2409 ( .A1(net31940), .A2(\u_div/CryTmp[7][18] ), .Y(n838) );
  NAND2X0_RVT U2410 ( .A1(\u_div/CryTmp[7][18] ), .A2(\u_div/PartRem[8][18] ), 
        .Y(n837) );
  IBUFFX4_RVT U2411 ( .A(net38347), .Y(net46859) );
  INVX1_RVT U2412 ( .A(net38347), .Y(net32518) );
  INVX1_RVT U2413 ( .A(net38347), .Y(net32520) );
  MUX21X1_RVT U2414 ( .A1(\u_div/PartRem[8][23] ), .A2(\u_div/SumTmp[7][23] ), 
        .S0(net46768), .Y(\u_div/PartRem[7][24] ) );
  INVX1_RVT U2415 ( .A(\u_div/SumTmp[7][22] ), .Y(net29680) );
  INVX0_RVT U2416 ( .A(\u_div/SumTmp[7][21] ), .Y(net29708) );
  NBUFFX4_RVT U2417 ( .A(n894), .Y(n883) );
  IBUFFX4_RVT U2418 ( .A(net48533), .Y(net52991) );
  INVX0_RVT U2419 ( .A(net52991), .Y(net52992) );
  INVX1_RVT U2420 ( .A(\u_div/PartRem[36][3] ), .Y(net52890) );
  MUX21X1_RVT U2421 ( .A1(net29837), .A2(net30696), .S0(net37570), .Y(net29846) );
  IBUFFX16_RVT U2422 ( .A(\u_div/SumTmp[13][7] ), .Y(net31196) );
  IBUFFX32_RVT U2423 ( .A(net42397), .Y(net42398) );
  NBUFFX8_RVT U2424 ( .A(net30992), .Y(net52536) );
  IBUFFX16_RVT U2425 ( .A(\u_div/SumTmp[30][2] ), .Y(net30992) );
  DELLN3X2_RVT U2426 ( .A(n240), .Y(net52520) );
  IBUFFX16_RVT U2427 ( .A(\u_div/SumTmp[12][11] ), .Y(net31155) );
  IBUFFX16_RVT U2428 ( .A(\u_div/CryTmp[6][18] ), .Y(n884) );
  INVX4_RVT U2429 ( .A(net29656), .Y(net51611) );
  IBUFFX16_RVT U2430 ( .A(\u_div/SumTmp[9][21] ), .Y(net29656) );
  IBUFFX32_RVT U2431 ( .A(net50339), .Y(net29821) );
  MUX21X2_RVT U2432 ( .A1(net29614), .A2(net30346), .S0(net40721), .Y(n1021)
         );
  IBUFFX16_RVT U2433 ( .A(\u_div/SumTmp[14][3] ), .Y(net30915) );
  IBUFFX4_RVT U2434 ( .A(n1055), .Y(\u_div/PartRem[38][6] ) );
  OR2X2_RVT U2435 ( .A1(\u_div/PartRem[7][24] ), .A2(\u_div/CryTmp[6][24] ), 
        .Y(net40656) );
  IBUFFX16_RVT U2436 ( .A(n1064), .Y(\u_div/PartRem[37][4] ) );
  IBUFFX16_RVT U2437 ( .A(\u_div/CryTmp[35][6] ), .Y(n1000) );
  IBUFFX16_RVT U2438 ( .A(n888), .Y(n886) );
  IBUFFX16_RVT U2439 ( .A(n886), .Y(n887) );
  IBUFFX4_RVT U2440 ( .A(net29841), .Y(\u_div/PartRem[36][8] ) );
  IBUFFX4_RVT U2441 ( .A(n1068), .Y(\u_div/PartRem[36][11] ) );
  IBUFFX4_RVT U2442 ( .A(n1070), .Y(\u_div/PartRem[35][12] ) );
  MUX21X1_RVT U2443 ( .A1(\u_div/SumTmp[38][2] ), .A2(\u_div/PartRem[39][2] ), 
        .S0(net46142), .Y(n964) );
  IBUFFX16_RVT U2444 ( .A(net37581), .Y(net46142) );
  IBUFFX16_RVT U2445 ( .A(\u_div/SumTmp[37][9] ), .Y(n1085) );
  MUX21X2_RVT U2446 ( .A1(n1029), .A2(n1040), .S0(net45257), .Y(net29685) );
  INVX4_RVT U2447 ( .A(net49213), .Y(net50185) );
  INVX2_RVT U2448 ( .A(net50185), .Y(net50186) );
  IBUFFX4_RVT U2449 ( .A(net49211), .Y(net50182) );
  IBUFFX4_RVT U2450 ( .A(net49211), .Y(net49213) );
  IBUFFX4_RVT U2451 ( .A(net49211), .Y(net49212) );
  IBUFFX16_RVT U2452 ( .A(n1059), .Y(\u_div/PartRem[37][9] ) );
  INVX8_RVT U2453 ( .A(n948), .Y(n889) );
  IBUFFX8_RVT U2454 ( .A(n889), .Y(n890) );
  INVX1_RVT U2455 ( .A(n1015), .Y(n985) );
  INVX1_RVT U2456 ( .A(\u_div/SumTmp[13][15] ), .Y(net31066) );
  INVX2_RVT U2457 ( .A(n929), .Y(n930) );
  IBUFFX16_RVT U2458 ( .A(n1071), .Y(\u_div/PartRem[35][11] ) );
  IBUFFX4_RVT U2459 ( .A(net49678), .Y(net49679) );
  INVX4_RVT U2460 ( .A(net30687), .Y(net49674) );
  IBUFFX4_RVT U2461 ( .A(net49674), .Y(net49675) );
  IBUFFX16_RVT U2462 ( .A(\u_div/SumTmp[27][11] ), .Y(net30687) );
  IBUFFX16_RVT U2463 ( .A(net29956), .Y(\u_div/PartRem[29][18] ) );
  IBUFFX16_RVT U2464 ( .A(\u_div/CryTmp[28][17] ), .Y(n891) );
  INVX4_RVT U2465 ( .A(n891), .Y(n892) );
  IBUFFX4_RVT U2466 ( .A(\u_div/SumTmp[27][12] ), .Y(net30639) );
  INVX4_RVT U2467 ( .A(n993), .Y(n893) );
  IBUFFX4_RVT U2468 ( .A(n893), .Y(n894) );
  INVX0_RVT U2469 ( .A(net49626), .Y(net49601) );
  INVX1_RVT U2470 ( .A(net29843), .Y(\u_div/PartRem[36][6] ) );
  IBUFFX4_RVT U2471 ( .A(n938), .Y(n1001) );
  IBUFFX16_RVT U2472 ( .A(b[22]), .Y(net31846) );
  NAND2X0_RVT U2473 ( .A1(net31800), .A2(\u_div/PartRem[2][23] ), .Y(n895) );
  NAND2X0_RVT U2474 ( .A1(n979), .A2(\u_div/PartRem[2][23] ), .Y(n896) );
  NAND2X0_RVT U2475 ( .A1(n979), .A2(net31800), .Y(n897) );
  NAND3X0_RVT U2476 ( .A1(n897), .A2(n896), .A3(n895), .Y(
        \u_div/CryTmp[1][24] ) );
  XOR3X1_RVT U2477 ( .A1(\u_div/PartRem[23][15] ), .A2(net32014), .A3(n214), 
        .Y(\u_div/SumTmp[22][15] ) );
  NAND2X0_RVT U2478 ( .A1(\u_div/PartRem[23][15] ), .A2(net32014), .Y(net49309) );
  NAND2X0_RVT U2479 ( .A1(net32014), .A2(n214), .Y(net49311) );
  XOR2X1_RVT U2480 ( .A1(n33), .A2(net31982), .Y(n898) );
  XOR2X2_RVT U2481 ( .A1(n898), .A2(\u_div/CryTmp[22][16] ), .Y(
        \u_div/SumTmp[22][16] ) );
  IBUFFX16_RVT U2482 ( .A(net29615), .Y(net49254) );
  IBUFFX4_RVT U2483 ( .A(net29821), .Y(\u_div/PartRem[38][9] ) );
  INVX2_RVT U2484 ( .A(net42938), .Y(net42939) );
  IBUFFX4_RVT U2485 ( .A(net47816), .Y(net49211) );
  IBUFFX32_RVT U2486 ( .A(\u_div/CryTmp[21][19] ), .Y(n899) );
  IBUFFX4_RVT U2487 ( .A(n899), .Y(n900) );
  IBUFFX4_RVT U2488 ( .A(n1066), .Y(\u_div/PartRem[36][9] ) );
  IBUFFX16_RVT U2489 ( .A(\u_div/CryTmp[27][13] ), .Y(n905) );
  INVX4_RVT U2490 ( .A(n905), .Y(n906) );
  INVX0_RVT U2491 ( .A(n907), .Y(n908) );
  INVX0_RVT U2492 ( .A(n909), .Y(n910) );
  IBUFFX16_RVT U2493 ( .A(net32542), .Y(net48339) );
  IBUFFX16_RVT U2494 ( .A(b[11]), .Y(net32130) );
  INVX0_RVT U2495 ( .A(n913), .Y(n914) );
  INVX0_RVT U2496 ( .A(n915), .Y(n916) );
  INVX0_RVT U2497 ( .A(n976), .Y(n977) );
  INVX0_RVT U2498 ( .A(n1172), .Y(\u_div/PartRem[2][10] ) );
  INVX1_RVT U2499 ( .A(net32624), .Y(net32620) );
  INVX1_RVT U2500 ( .A(net47709), .Y(net32624) );
  MUX21X1_RVT U2501 ( .A1(\u_div/PartRem[23][23] ), .A2(\u_div/SumTmp[22][23] ), .S0(net32610), .Y(\u_div/PartRem[22][24] ) );
  INVX4_RVT U2502 ( .A(net46241), .Y(net48758) );
  IBUFFX16_RVT U2503 ( .A(net48758), .Y(net48759) );
  IBUFFX16_RVT U2504 ( .A(net31261), .Y(net43884) );
  INVX1_RVT U2505 ( .A(\u_div/PartRem[3][8] ), .Y(n935) );
  IBUFFX32_RVT U2506 ( .A(\u_div/CryTmp[35][9] ), .Y(n927) );
  INVX1_RVT U2507 ( .A(n927), .Y(n928) );
  IBUFFX16_RVT U2508 ( .A(net47688), .Y(net48670) );
  INVX4_RVT U2509 ( .A(net48670), .Y(net48671) );
  NOR2X4_RVT U2510 ( .A1(\u_div/CryTmp[13][24] ), .A2(\u_div/PartRem[14][24] ), 
        .Y(net47688) );
  IBUFFX16_RVT U2511 ( .A(net39869), .Y(net39872) );
  INVX1_RVT U2512 ( .A(net48638), .Y(net48639) );
  INVX1_RVT U2513 ( .A(net29899), .Y(\u_div/PartRem[32][15] ) );
  IBUFFX16_RVT U2514 ( .A(\u_div/CryTmp[6][21] ), .Y(n929) );
  INVX2_RVT U2515 ( .A(n883), .Y(n994) );
  INVX1_RVT U2516 ( .A(net29658), .Y(\u_div/PartRem[7][21] ) );
  INVX1_RVT U2517 ( .A(n1029), .Y(\u_div/PartRem[7][20] ) );
  INVX1_RVT U2518 ( .A(net29661), .Y(\u_div/PartRem[7][19] ) );
  IBUFFX16_RVT U2519 ( .A(n981), .Y(n947) );
  IBUFFX16_RVT U2520 ( .A(n989), .Y(n990) );
  IBUFFX16_RVT U2521 ( .A(\u_div/CryTmp[33][13] ), .Y(n931) );
  INVX4_RVT U2522 ( .A(n931), .Y(n932) );
  INVX1_RVT U2523 ( .A(\u_div/CryTmp[28][16] ), .Y(n933) );
  IBUFFX4_RVT U2524 ( .A(n933), .Y(n934) );
  INVX1_RVT U2525 ( .A(n1194), .Y(\u_div/PartRem[14][23] ) );
  IBUFFX4_RVT U2526 ( .A(net48384), .Y(net48385) );
  INVX1_RVT U2527 ( .A(net48339), .Y(net48340) );
  INVX1_RVT U2528 ( .A(net48339), .Y(net48341) );
  INVX1_RVT U2529 ( .A(net48339), .Y(net48342) );
  INVX1_RVT U2530 ( .A(n1045), .Y(\u_div/PartRem[3][18] ) );
  INVX0_RVT U2531 ( .A(n1004), .Y(n1005) );
  INVX1_RVT U2532 ( .A(n1046), .Y(\u_div/PartRem[3][17] ) );
  INVX1_RVT U2533 ( .A(n1044), .Y(\u_div/PartRem[3][19] ) );
  INVX2_RVT U2534 ( .A(n1000), .Y(n937) );
  INVX1_RVT U2535 ( .A(n996), .Y(n997) );
  INVX0_RVT U2536 ( .A(n954), .Y(n955) );
  IBUFFX4_RVT U2537 ( .A(\u_div/CryTmp[37][8] ), .Y(n939) );
  INVX1_RVT U2538 ( .A(n939), .Y(n940) );
  IBUFFX16_RVT U2539 ( .A(\u_div/CryTmp[7][16] ), .Y(n943) );
  INVX2_RVT U2540 ( .A(n991), .Y(n992) );
  INVX0_RVT U2541 ( .A(n965), .Y(n966) );
  IBUFFX4_RVT U2542 ( .A(net47978), .Y(net47979) );
  INVX1_RVT U2543 ( .A(n1042), .Y(\u_div/PartRem[3][21] ) );
  INVX0_RVT U2544 ( .A(net29801), .Y(\u_div/PartRem[3][20] ) );
  IBUFFX32_RVT U2545 ( .A(n947), .Y(n948) );
  NBUFFX2_RVT U2546 ( .A(net42515), .Y(net45587) );
  INVX1_RVT U2547 ( .A(net45669), .Y(net45677) );
  INVX1_RVT U2548 ( .A(net42548), .Y(net42512) );
  NBUFFX2_RVT U2549 ( .A(net42512), .Y(net45588) );
  INVX1_RVT U2550 ( .A(b[18]), .Y(net31952) );
  NOR4X1_RVT U2551 ( .A1(net31255), .A2(n1229), .A3(net32210), .A4(n121), .Y(
        net47816) );
  INVX1_RVT U2552 ( .A(net32156), .Y(net32154) );
  INVX1_RVT U2553 ( .A(n952), .Y(n953) );
  INVX1_RVT U2554 ( .A(n890), .Y(quotient[2]) );
  INVX1_RVT U2555 ( .A(net46961), .Y(net46962) );
  INVX1_RVT U2556 ( .A(net44967), .Y(net46961) );
  OR2X1_RVT U2557 ( .A1(\u_div/PartRem[15][24] ), .A2(\u_div/CryTmp[14][24] ), 
        .Y(net47718) );
  INVX1_RVT U2558 ( .A(b[16]), .Y(net32002) );
  INVX1_RVT U2559 ( .A(n1016), .Y(n983) );
  INVX1_RVT U2560 ( .A(n1007), .Y(n1016) );
  INVX1_RVT U2561 ( .A(n983), .Y(quotient[1]) );
  INVX1_RVT U2562 ( .A(\u_div/SumTmp[24][2] ), .Y(net31116) );
  INVX1_RVT U2563 ( .A(\u_div/SumTmp[24][1] ), .Y(net31134) );
  INVX1_RVT U2564 ( .A(b[15]), .Y(net32032) );
  AND3X1_RVT U2565 ( .A1(net31952), .A2(net32386), .A3(net31930), .Y(n949) );
  XNOR2X1_RVT U2566 ( .A1(\u_div/CryTmp[7][18] ), .A2(n1002), .Y(n950) );
  INVX0_RVT U2567 ( .A(net45669), .Y(net45671) );
  INVX1_RVT U2568 ( .A(b[19]), .Y(net31930) );
  INVX1_RVT U2569 ( .A(\u_div/SumTmp[26][7] ), .Y(net30962) );
  INVX1_RVT U2570 ( .A(\u_div/SumTmp[33][11] ), .Y(net30210) );
  INVX1_RVT U2571 ( .A(net47979), .Y(net44967) );
  INVX0_RVT U2572 ( .A(\u_div/PartRem[2][24] ), .Y(n974) );
  OR2X1_RVT U2573 ( .A1(\u_div/PartRem[10][24] ), .A2(\u_div/CryTmp[9][24] ), 
        .Y(net46550) );
  IBUFFX16_RVT U2574 ( .A(\u_div/SumTmp[13][13] ), .Y(net31105) );
  MUX21X1_RVT U2575 ( .A1(net29854), .A2(net30598), .S0(net37563), .Y(net46421) );
  IBUFFX16_RVT U2576 ( .A(\u_div/SumTmp[13][11] ), .Y(net31140) );
  IBUFFX16_RVT U2577 ( .A(\u_div/SumTmp[8][22] ), .Y(net29654) );
  IBUFFX4_RVT U2578 ( .A(net48759), .Y(net46242) );
  IBUFFX16_RVT U2579 ( .A(\u_div/SumTmp[35][8] ), .Y(net30260) );
  IBUFFX4_RVT U2580 ( .A(\u_div/CryTmp[9][23] ), .Y(n967) );
  IBUFFX16_RVT U2581 ( .A(\u_div/PartRem[1][16] ), .Y(n969) );
  IBUFFX16_RVT U2582 ( .A(n1067), .Y(\u_div/PartRem[36][7] ) );
  IBUFFX16_RVT U2583 ( .A(\u_div/PartRem[1][15] ), .Y(n971) );
  MUX21X1_RVT U2584 ( .A1(net31530), .A2(n1012), .S0(n171), .Y(net29820) );
  NAND2X0_RVT U2585 ( .A1(n974), .A2(n975), .Y(n973) );
  IBUFFX16_RVT U2586 ( .A(n973), .Y(n1007) );
  IBUFFX8_RVT U2587 ( .A(\u_div/CryTmp[1][24] ), .Y(n975) );
  IBUFFX16_RVT U2588 ( .A(\u_div/SumTmp[28][11] ), .Y(n1186) );
  IBUFFX16_RVT U2589 ( .A(\u_div/SumTmp[14][9] ), .Y(net31157) );
  INVX1_RVT U2590 ( .A(\u_div/SumTmp[8][18] ), .Y(net29796) );
  IBUFFX4_RVT U2591 ( .A(net45669), .Y(net45678) );
  NOR2X1_RVT U2592 ( .A1(net31255), .A2(n1223), .Y(net37556) );
  INVX0_RVT U2593 ( .A(net42548), .Y(net45599) );
  INVX0_RVT U2594 ( .A(net42548), .Y(net45601) );
  INVX0_RVT U2595 ( .A(net42548), .Y(net45602) );
  INVX0_RVT U2596 ( .A(net42548), .Y(net45603) );
  INVX0_RVT U2597 ( .A(net42548), .Y(net45604) );
  IBUFFX16_RVT U2598 ( .A(\u_div/SumTmp[15][7] ), .Y(net31173) );
  INVX1_RVT U2599 ( .A(\u_div/SumTmp[9][2] ), .Y(net30468) );
  IBUFFX4_RVT U2600 ( .A(net46550), .Y(net45541) );
  IBUFFX16_RVT U2601 ( .A(\u_div/SumTmp[8][3] ), .Y(net30466) );
  NOR2X1_RVT U2602 ( .A1(\u_div/CryTmp[2][24] ), .A2(\u_div/PartRem[3][24] ), 
        .Y(n1008) );
  IBUFFX16_RVT U2603 ( .A(\u_div/SumTmp[25][4] ), .Y(net31056) );
  INVX2_RVT U2604 ( .A(net29755), .Y(\u_div/PartRem[46][1] ) );
  IBUFFX16_RVT U2605 ( .A(\u_div/SumTmp[24][8] ), .Y(net30986) );
  INVX8_RVT U2606 ( .A(n1102), .Y(\u_div/PartRem[23][11] ) );
  IBUFFX16_RVT U2607 ( .A(\u_div/SumTmp[24][9] ), .Y(net30960) );
  MUX21X1_RVT U2608 ( .A1(net30022), .A2(net30733), .S0(quotient[25]), .Y(
        net45295) );
  NOR2X1_RVT U2609 ( .A1(\u_div/PartRem[21][24] ), .A2(\u_div/CryTmp[20][24] ), 
        .Y(net38343) );
  MUX21X1_RVT U2610 ( .A1(net30801), .A2(n75), .S0(quotient[12]), .Y(net45288)
         );
  INVX2_RVT U2611 ( .A(n95), .Y(n1114) );
  IBUFFX16_RVT U2612 ( .A(\u_div/SumTmp[12][15] ), .Y(net31085) );
  IBUFFX16_RVT U2613 ( .A(\u_div/SumTmp[12][14] ), .Y(net31104) );
  IBUFFX16_RVT U2614 ( .A(\u_div/SumTmp[14][6] ), .Y(net31197) );
  IBUFFX16_RVT U2615 ( .A(\u_div/SumTmp[12][19] ), .Y(net30998) );
  IBUFFX16_RVT U2616 ( .A(\u_div/SumTmp[12][20] ), .Y(net30974) );
  IBUFFX16_RVT U2617 ( .A(\u_div/SumTmp[13][9] ), .Y(net31171) );
  IBUFFX16_RVT U2618 ( .A(\u_div/SumTmp[27][3] ), .Y(net31036) );
  INVX1_RVT U2619 ( .A(net47979), .Y(net45007) );
  MUX21X1_RVT U2620 ( .A1(net30758), .A2(net31123), .S0(net32554), .Y(net45002) );
  IBUFFX16_RVT U2621 ( .A(\u_div/SumTmp[14][11] ), .Y(net31124) );
  IBUFFX16_RVT U2622 ( .A(\u_div/SumTmp[14][8] ), .Y(net31172) );
  MUX21X1_RVT U2623 ( .A1(net29752), .A2(net30421), .S0(net45594), .Y(n1050)
         );
  MUX21X1_RVT U2624 ( .A1(net29818), .A2(net30554), .S0(net37581), .Y(n1057)
         );
  IBUFFX4_RVT U2625 ( .A(\u_div/SumTmp[17][17] ), .Y(net30869) );
  IBUFFX16_RVT U2626 ( .A(\u_div/SumTmp[17][18] ), .Y(net30821) );
  IBUFFX4_RVT U2627 ( .A(\u_div/CryTmp[28][18] ), .Y(n989) );
  IBUFFX16_RVT U2628 ( .A(\u_div/SumTmp[29][14] ), .Y(net30254) );
  IBUFFX16_RVT U2629 ( .A(\u_div/SumTmp[35][5] ), .Y(net30599) );
  IBUFFX16_RVT U2630 ( .A(\u_div/SumTmp[24][4] ), .Y(net31077) );
  IBUFFX16_RVT U2631 ( .A(\u_div/SumTmp[13][17] ), .Y(net31022) );
  IBUFFX2_RVT U2632 ( .A(\u_div/PartRem[38][9] ), .Y(net44466) );
  IBUFFX16_RVT U2633 ( .A(net29822), .Y(\u_div/PartRem[38][8] ) );
  IBUFFX16_RVT U2634 ( .A(n1054), .Y(\u_div/PartRem[38][7] ) );
  MUX21X2_RVT U2635 ( .A1(n1055), .A2(n1128), .S0(net37242), .Y(n1061) );
  IBUFFX16_RVT U2636 ( .A(n1056), .Y(\u_div/PartRem[38][5] ) );
  IBUFFX16_RVT U2637 ( .A(n1057), .Y(\u_div/PartRem[38][4] ) );
  IBUFFX16_RVT U2638 ( .A(n1060), .Y(\u_div/PartRem[37][8] ) );
  IBUFFX16_RVT U2639 ( .A(n1061), .Y(\u_div/PartRem[37][7] ) );
  IBUFFX16_RVT U2640 ( .A(\u_div/CryTmp[36][7] ), .Y(n991) );
  IBUFFX4_RVT U2641 ( .A(\u_div/SumTmp[35][11] ), .Y(n1083) );
  IBUFFX16_RVT U2642 ( .A(\u_div/CryTmp[27][19] ), .Y(n993) );
  MUX21X1_RVT U2643 ( .A1(net29698), .A2(net46608), .S0(net50726), .Y(n995) );
  IBUFFX4_RVT U2644 ( .A(n1193), .Y(\u_div/PartRem[14][22] ) );
  IBUFFX4_RVT U2645 ( .A(net30748), .Y(\u_div/PartRem[14][21] ) );
  MUX21X2_RVT U2646 ( .A1(n1013), .A2(n1017), .S0(n1086), .Y(net29755) );
  IBUFFX4_RVT U2647 ( .A(\u_div/CryTmp[34][11] ), .Y(net44063) );
  INVX2_RVT U2648 ( .A(net44063), .Y(net44064) );
  INVX1_RVT U2649 ( .A(net43884), .Y(net43885) );
  IBUFFX4_RVT U2650 ( .A(n1069), .Y(\u_div/PartRem[36][10] ) );
  IBUFFX16_RVT U2651 ( .A(net31255), .Y(net43354) );
  NAND2X0_RVT U2652 ( .A1(\u_div/CryTmp[37][10] ), .A2(net43354), .Y(net43355)
         );
  IBUFFX16_RVT U2653 ( .A(\u_div/SumTmp[35][9] ), .Y(n1122) );
  IBUFFX16_RVT U2654 ( .A(\u_div/SumTmp[31][11] ), .Y(net30499) );
  MUX21X1_RVT U2655 ( .A1(net29731), .A2(net30304), .S0(net45581), .Y(n1036)
         );
  IBUFFX4_RVT U2656 ( .A(\u_div/CryTmp[31][15] ), .Y(net42397) );
  IBUFFX16_RVT U2657 ( .A(net32592), .Y(net42365) );
  IBUFFX16_RVT U2658 ( .A(net47718), .Y(net42357) );
  IBUFFX4_RVT U2659 ( .A(net30182), .Y(\u_div/PartRem[22][17] ) );
  IBUFFX16_RVT U2660 ( .A(net30178), .Y(\u_div/PartRem[22][20] ) );
  AND3X1_RVT U2661 ( .A1(net32032), .A2(net31974), .A3(net32002), .Y(n1095) );
  INVX2_RVT U2662 ( .A(b[17]), .Y(net31974) );
  XNOR2X1_RVT U2663 ( .A1(a[25]), .A2(net32406), .Y(net41046) );
  MUX21X1_RVT U2664 ( .A1(\u_div/SumTmp[8][10] ), .A2(\u_div/PartRem[9][10] ), 
        .S0(net40717), .Y(n1003) );
  IBUFFX16_RVT U2665 ( .A(net47729), .Y(net40724) );
  INVX0_RVT U2666 ( .A(net29662), .Y(\u_div/PartRem[7][18] ) );
  IBUFFX4_RVT U2667 ( .A(net40724), .Y(net40717) );
  INVX2_RVT U2668 ( .A(net39872), .Y(net39874) );
  AND2X1_RVT U2669 ( .A1(net39870), .A2(\u_div/CryTmp[31][16] ), .Y(net39869)
         );
  NOR2X1_RVT U2670 ( .A1(net32104), .A2(net31287), .Y(n1006) );
  INVX0_RVT U2671 ( .A(\u_div/CryTmp[11][1] ), .Y(\u_div/SumTmp[7][0] ) );
  INVX0_RVT U2672 ( .A(\u_div/CryTmp[11][1] ), .Y(\u_div/SumTmp[6][0] ) );
  INVX0_RVT U2673 ( .A(\u_div/CryTmp[11][1] ), .Y(\u_div/SumTmp[9][0] ) );
  INVX0_RVT U2674 ( .A(net30293), .Y(\*cell*33726/net34245 ) );
  INVX0_RVT U2675 ( .A(\u_div/CryTmp[11][1] ), .Y(\u_div/SumTmp[11][0] ) );
  INVX0_RVT U2676 ( .A(net30945), .Y(\*cell*33681/net34095 ) );
  INVX0_RVT U2677 ( .A(\u_div/CryTmp[11][1] ), .Y(\u_div/SumTmp[8][0] ) );
  INVX0_RVT U2678 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[12][0] ) );
  INVX0_RVT U2679 ( .A(net30943), .Y(\*cell*33684/net34105 ) );
  INVX0_RVT U2680 ( .A(\u_div/CryTmp[11][1] ), .Y(\u_div/SumTmp[5][0] ) );
  INVX0_RVT U2681 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[18][0] ) );
  INVX0_RVT U2682 ( .A(net30910), .Y(\*cell*33702/net34165 ) );
  INVX0_RVT U2683 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[15][0] ) );
  INVX0_RVT U2684 ( .A(net30931), .Y(\*cell*33693/net34135 ) );
  INVX0_RVT U2685 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[14][0] ) );
  INVX0_RVT U2686 ( .A(net30936), .Y(\*cell*33690/net34125 ) );
  INVX0_RVT U2687 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[13][0] ) );
  INVX0_RVT U2688 ( .A(net30940), .Y(\*cell*33687/net34115 ) );
  INVX0_RVT U2689 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[16][0] ) );
  INVX0_RVT U2690 ( .A(net30925), .Y(\*cell*33696/net34145 ) );
  INVX0_RVT U2691 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[20][0] ) );
  INVX0_RVT U2692 ( .A(net31203), .Y(\*cell*33669/net34055 ) );
  INVX0_RVT U2693 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[21][0] ) );
  INVX0_RVT U2694 ( .A(net31192), .Y(\*cell*33672/net34065 ) );
  INVX0_RVT U2695 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[19][0] ) );
  INVX0_RVT U2696 ( .A(net31213), .Y(\*cell*33666/net34045 ) );
  INVX0_RVT U2697 ( .A(\u_div/CryTmp[22][1] ), .Y(\u_div/SumTmp[22][0] ) );
  INVX0_RVT U2698 ( .A(net31180), .Y(\*cell*33675/net34075 ) );
  INVX1_RVT U2699 ( .A(n1135), .Y(\u_div/PartRem[2][4] ) );
  INVX1_RVT U2700 ( .A(\u_div/SumTmp[2][3] ), .Y(n1136) );
  INVX1_RVT U2701 ( .A(n1131), .Y(\u_div/PartRem[2][6] ) );
  INVX1_RVT U2702 ( .A(\u_div/SumTmp[2][5] ), .Y(n1132) );
  INVX1_RVT U2703 ( .A(n1129), .Y(\u_div/PartRem[2][7] ) );
  INVX1_RVT U2704 ( .A(\u_div/SumTmp[2][6] ), .Y(n1130) );
  INVX1_RVT U2705 ( .A(n1191), .Y(\u_div/PartRem[15][23] ) );
  INVX1_RVT U2706 ( .A(\u_div/SumTmp[13][22] ), .Y(n1197) );
  INVX1_RVT U2707 ( .A(\u_div/SumTmp[12][22] ), .Y(net30864) );
  INVX1_RVT U2708 ( .A(n1202), .Y(\u_div/PartRem[10][23] ) );
  INVX1_RVT U2709 ( .A(\u_div/SumTmp[9][22] ), .Y(n1020) );
  INVX1_RVT U2710 ( .A(n1030), .Y(\u_div/PartRem[7][23] ) );
  INVX1_RVT U2711 ( .A(n1150), .Y(\u_div/PartRem[2][20] ) );
  INVX1_RVT U2712 ( .A(\u_div/SumTmp[2][19] ), .Y(n1151) );
  INVX1_RVT U2713 ( .A(n1147), .Y(\u_div/PartRem[2][21] ) );
  INVX1_RVT U2714 ( .A(\u_div/SumTmp[2][20] ), .Y(n1148) );
  INVX1_RVT U2715 ( .A(n1144), .Y(\u_div/PartRem[2][22] ) );
  INVX1_RVT U2716 ( .A(\u_div/SumTmp[2][21] ), .Y(n1145) );
  INVX1_RVT U2717 ( .A(net30180), .Y(\u_div/PartRem[22][19] ) );
  INVX1_RVT U2718 ( .A(net29981), .Y(\u_div/PartRem[28][12] ) );
  INVX1_RVT U2719 ( .A(net29978), .Y(\u_div/PartRem[28][15] ) );
  INVX1_RVT U2720 ( .A(n1075), .Y(\u_div/PartRem[29][15] ) );
  INVX1_RVT U2721 ( .A(net29682), .Y(\u_div/PartRem[10][20] ) );
  INVX1_RVT U2722 ( .A(net30702), .Y(\u_div/PartRem[15][20] ) );
  INVX1_RVT U2723 ( .A(n1189), .Y(\u_div/PartRem[15][22] ) );
  INVX1_RVT U2724 ( .A(net29844), .Y(\u_div/PartRem[36][5] ) );
  INVX1_RVT U2725 ( .A(n1190), .Y(\u_div/PartRem[15][21] ) );
  INVX1_RVT U2726 ( .A(n1022), .Y(\u_div/PartRem[8][15] ) );
  INVX1_RVT U2727 ( .A(net29665), .Y(\u_div/PartRem[7][15] ) );
  INVX1_RVT U2728 ( .A(net29710), .Y(\u_div/PartRem[10][19] ) );
  INVX1_RVT U2729 ( .A(net29655), .Y(\u_div/PartRem[10][21] ) );
  INVX1_RVT U2730 ( .A(n1137), .Y(\u_div/PartRem[2][3] ) );
  INVX1_RVT U2731 ( .A(\u_div/SumTmp[2][2] ), .Y(n1138) );
  INVX1_RVT U2732 ( .A(n1133), .Y(\u_div/PartRem[2][5] ) );
  INVX1_RVT U2733 ( .A(\u_div/SumTmp[2][4] ), .Y(n1134) );
  INVX1_RVT U2734 ( .A(\u_div/SumTmp[2][8] ), .Y(n1175) );
  INVX1_RVT U2735 ( .A(n1062), .Y(\u_div/PartRem[37][6] ) );
  INVX1_RVT U2736 ( .A(n1099), .Y(\u_div/PartRem[23][14] ) );
  INVX1_RVT U2737 ( .A(net29982), .Y(\u_div/PartRem[28][11] ) );
  INVX1_RVT U2738 ( .A(net29979), .Y(\u_div/PartRem[28][14] ) );
  INVX1_RVT U2739 ( .A(net30033), .Y(\u_div/PartRem[25][22] ) );
  INVX1_RVT U2740 ( .A(n1080), .Y(\u_div/PartRem[29][10] ) );
  INVX1_RVT U2741 ( .A(n1079), .Y(\u_div/PartRem[29][11] ) );
  INVX1_RVT U2742 ( .A(n1076), .Y(\u_div/PartRem[29][14] ) );
  INVX1_RVT U2743 ( .A(net29666), .Y(\u_div/PartRem[7][14] ) );
  INVX1_RVT U2744 ( .A(n1049), .Y(\u_div/PartRem[3][14] ) );
  INVX1_RVT U2745 ( .A(net29637), .Y(\u_div/PartRem[8][17] ) );
  INVX1_RVT U2746 ( .A(net29663), .Y(\u_div/PartRem[7][17] ) );
  INVX1_RVT U2747 ( .A(net30185), .Y(\u_div/PartRem[22][14] ) );
  INVX1_RVT U2748 ( .A(net29669), .Y(\u_div/PartRem[7][11] ) );
  INVX1_RVT U2749 ( .A(net29874), .Y(\u_div/PartRem[34][11] ) );
  INVX1_RVT U2750 ( .A(net30186), .Y(\u_div/PartRem[22][13] ) );
  INVX1_RVT U2751 ( .A(net29667), .Y(\u_div/PartRem[7][13] ) );
  INVX1_RVT U2752 ( .A(n1050), .Y(\u_div/PartRem[3][13] ) );
  INVX1_RVT U2753 ( .A(n1139), .Y(\u_div/PartRem[2][2] ) );
  INVX1_RVT U2754 ( .A(\u_div/SumTmp[2][1] ), .Y(n1140) );
  NOR2X0_RVT U2755 ( .A1(\u_div/CryTmp[12][24] ), .A2(\u_div/PartRem[13][24] ), 
        .Y(net38337) );
  INVX1_RVT U2756 ( .A(n1170), .Y(\u_div/PartRem[2][13] ) );
  INVX1_RVT U2757 ( .A(n1162), .Y(\u_div/PartRem[2][16] ) );
  INVX1_RVT U2758 ( .A(n1159), .Y(\u_div/PartRem[2][17] ) );
  MUX21X1_RVT U2759 ( .A1(\u_div/PartRem[7][22] ), .A2(\u_div/SumTmp[6][22] ), 
        .S0(net45257), .Y(n1009) );
  INVX1_RVT U2760 ( .A(net30184), .Y(\u_div/PartRem[22][15] ) );
  INVX1_RVT U2761 ( .A(n1038), .Y(\u_div/PartRem[3][3] ) );
  INVX1_RVT U2762 ( .A(net30183), .Y(\u_div/PartRem[22][16] ) );
  INVX1_RVT U2763 ( .A(n1047), .Y(\u_div/PartRem[3][16] ) );
  INVX1_RVT U2764 ( .A(n1101), .Y(\u_div/PartRem[23][12] ) );
  INVX1_RVT U2765 ( .A(n1018), .Y(\u_div/PartRem[8][9] ) );
  INVX1_RVT U2766 ( .A(net29873), .Y(\u_div/PartRem[34][12] ) );
  INVX1_RVT U2767 ( .A(n1063), .Y(\u_div/PartRem[37][5] ) );
  INVX1_RVT U2768 ( .A(n1078), .Y(\u_div/PartRem[29][12] ) );
  NAND2X0_RVT U2769 ( .A1(net47690), .A2(\u_div/CryTmp[28][19] ), .Y(net31310)
         );
  MUX21X1_RVT U2770 ( .A1(n1011), .A2(\u_div/SumTmp[2][11] ), .S0(n987), .Y(
        n1010) );
  INVX1_RVT U2771 ( .A(n1165), .Y(\u_div/PartRem[2][15] ) );
  INVX1_RVT U2772 ( .A(n1156), .Y(\u_div/PartRem[2][18] ) );
  INVX1_RVT U2773 ( .A(net31276), .Y(net31272) );
  INVX1_RVT U2774 ( .A(n1037), .Y(\u_div/PartRem[3][4] ) );
  INVX1_RVT U2775 ( .A(n1039), .Y(\u_div/PartRem[3][2] ) );
  INVX1_RVT U2776 ( .A(n1100), .Y(\u_div/PartRem[23][13] ) );
  INVX1_RVT U2777 ( .A(net30130), .Y(\u_div/PartRem[23][10] ) );
  INVX1_RVT U2778 ( .A(n1027), .Y(\u_div/PartRem[8][10] ) );
  INVX1_RVT U2779 ( .A(net29670), .Y(\u_div/PartRem[7][10] ) );
  INVX1_RVT U2780 ( .A(n1077), .Y(\u_div/PartRem[29][13] ) );
  AND2X1_RVT U2781 ( .A1(net32092), .A2(net32068), .Y(net31250) );
  AND2X1_RVT U2782 ( .A1(net31964), .A2(net31952), .Y(n1222) );
  INVX1_RVT U2783 ( .A(n1141), .Y(\u_div/PartRem[2][1] ) );
  MUX21X1_RVT U2784 ( .A1(\u_div/PartRem[2][10] ), .A2(\u_div/SumTmp[1][10] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][11] ) );
  INVX1_RVT U2785 ( .A(net30314), .Y(\*cell*33717/net34215 ) );
  INVX1_RVT U2786 ( .A(net30308), .Y(\*cell*33720/net34225 ) );
  INVX1_RVT U2787 ( .A(net30301), .Y(\*cell*33723/net34235 ) );
  INVX1_RVT U2788 ( .A(n1043), .Y(\u_div/PartRem[3][1] ) );
  XOR2X1_RVT U2789 ( .A1(a[28]), .A2(net32406), .Y(net37263) );
  XOR2X1_RVT U2790 ( .A1(a[30]), .A2(net32406), .Y(net37261) );
  XOR2X1_RVT U2791 ( .A1(a[39]), .A2(net32408), .Y(n1012) );
  XOR2X1_RVT U2792 ( .A1(a[41]), .A2(net32408), .Y(net37256) );
  XOR2X1_RVT U2793 ( .A1(a[32]), .A2(net32406), .Y(net37254) );
  XOR2X1_RVT U2794 ( .A1(a[26]), .A2(net32406), .Y(net37253) );
  XOR2X1_RVT U2795 ( .A1(a[40]), .A2(net32408), .Y(net37252) );
  XOR2X1_RVT U2796 ( .A1(a[36]), .A2(net32408), .Y(net37251) );
  XOR2X1_RVT U2797 ( .A1(a[37]), .A2(net32408), .Y(net37249) );
  XOR2X1_RVT U2798 ( .A1(a[27]), .A2(net32406), .Y(net37248) );
  XOR2X1_RVT U2799 ( .A1(a[35]), .A2(net32406), .Y(net37247) );
  XOR2X1_RVT U2800 ( .A1(a[34]), .A2(net32406), .Y(net37246) );
  XOR2X1_RVT U2801 ( .A1(a[31]), .A2(net32406), .Y(net37244) );
  INVX1_RVT U2802 ( .A(a[41]), .Y(net31498) );
  INVX1_RVT U2803 ( .A(net32106), .Y(net32104) );
  XOR2X1_RVT U2804 ( .A1(a[33]), .A2(net32406), .Y(net37231) );
  XOR2X1_RVT U2805 ( .A1(a[24]), .A2(net32406), .Y(net37229) );
  XOR2X1_RVT U2806 ( .A1(a[23]), .A2(\u_div/CryTmp[22][1] ), .Y(net37228) );
  OR2X1_RVT U2807 ( .A1(net32408), .A2(a[45]), .Y(\u_div/CryTmp[45][1] ) );
  XOR2X1_RVT U2808 ( .A1(a[43]), .A2(net32408), .Y(net37224) );
  XOR2X1_RVT U2809 ( .A1(a[46]), .A2(net32408), .Y(n1013) );
  OR2X1_RVT U2810 ( .A1(n1108), .A2(n1109), .Y(net37219) );
  XOR2X1_RVT U2811 ( .A1(a[45]), .A2(net32408), .Y(net37220) );
  NOR2X0_RVT U2812 ( .A1(net32408), .A2(a[46]), .Y(n1014) );
  INVX1_RVT U2813 ( .A(a[40]), .Y(net31514) );
  INVX1_RVT U2814 ( .A(a[45]), .Y(net31434) );
  INVX1_RVT U2815 ( .A(b[23]), .Y(net31822) );
  INVX1_RVT U2816 ( .A(a[46]), .Y(n1017) );
  XOR2X1_RVT U2817 ( .A1(a[42]), .A2(net32408), .Y(net37184) );
  INVX1_RVT U2818 ( .A(a[42]), .Y(net31482) );
  INVX1_RVT U2819 ( .A(a[43]), .Y(net31466) );
  INVX1_RVT U2820 ( .A(a[39]), .Y(net31530) );
  INVX1_RVT U2821 ( .A(a[37]), .Y(net31562) );
  INVX1_RVT U2822 ( .A(a[36]), .Y(net31578) );
  INVX1_RVT U2823 ( .A(a[35]), .Y(net31594) );
  INVX1_RVT U2824 ( .A(a[34]), .Y(net31610) );
  INVX1_RVT U2825 ( .A(a[33]), .Y(net31626) );
  INVX1_RVT U2826 ( .A(a[32]), .Y(net31642) );
  INVX1_RVT U2827 ( .A(a[31]), .Y(net31658) );
  AND2X1_RVT U2828 ( .A1(quotient[1]), .A2(\u_div/SumTmp[5][0] ), .Y(
        \u_div/PartRem[1][1] ) );
  INVX1_RVT U2829 ( .A(a[30]), .Y(net31674) );
  INVX1_RVT U2830 ( .A(a[28]), .Y(net31706) );
  INVX1_RVT U2831 ( .A(a[27]), .Y(net31722) );
  INVX1_RVT U2832 ( .A(a[26]), .Y(net31738) );
  INVX1_RVT U2833 ( .A(a[24]), .Y(net31770) );
  INVX1_RVT U2834 ( .A(a[23]), .Y(net31786) );
  INVX1_RVT U2835 ( .A(b[12]), .Y(net32106) );
  INVX1_RVT U2836 ( .A(b[21]), .Y(net31874) );
  INVX1_RVT U2837 ( .A(b[20]), .Y(net31902) );
  NAND2X0_RVT U2838 ( .A1(n987), .A2(\u_div/SumTmp[5][0] ), .Y(n1141) );
  INVX1_RVT U2839 ( .A(n1074), .Y(\u_div/PartRem[29][16] ) );
  INVX1_RVT U2840 ( .A(n1153), .Y(\u_div/PartRem[2][19] ) );
  MUX21X1_RVT U2841 ( .A1(\u_div/PartRem[10][23] ), .A2(\u_div/SumTmp[9][23] ), 
        .S0(net32530), .Y(\u_div/PartRem[9][24] ) );
  MUX21X1_RVT U2842 ( .A1(net29606), .A2(net29654), .S0(net40718), .Y(net29653) );
  MUX21X1_RVT U2843 ( .A1(\u_div/PartRem[7][23] ), .A2(\u_div/SumTmp[6][23] ), 
        .S0(net45257), .Y(\u_div/PartRem[6][24] ) );
  MUX21X1_RVT U2844 ( .A1(net29631), .A2(net29680), .S0(net46859), .Y(n1030)
         );
  INVX0_RVT U2845 ( .A(\u_div/SumTmp[9][20] ), .Y(net29683) );
  MUX21X1_RVT U2846 ( .A1(n1009), .A2(\u_div/SumTmp[5][23] ), .S0(net44755), 
        .Y(\u_div/PartRem[5][24] ) );
  MUX21X1_RVT U2847 ( .A1(net29632), .A2(net29708), .S0(net46768), .Y(n1028)
         );
  INVX0_RVT U2848 ( .A(\u_div/SumTmp[8][20] ), .Y(net29709) );
  INVX0_RVT U2849 ( .A(\u_div/SumTmp[9][19] ), .Y(net29711) );
  MUX21X1_RVT U2850 ( .A1(net29658), .A2(n1031), .S0(net45257), .Y(net29684)
         );
  INVX0_RVT U2851 ( .A(\u_div/SumTmp[6][21] ), .Y(n1031) );
  INVX0_RVT U2852 ( .A(\u_div/SumTmp[6][20] ), .Y(n1040) );
  MUX21X1_RVT U2853 ( .A1(net29635), .A2(net29795), .S0(net46859), .Y(n1029)
         );
  INVX0_RVT U2854 ( .A(\u_div/SumTmp[7][19] ), .Y(net29795) );
  MUX21X1_RVT U2855 ( .A1(\u_div/PartRem[3][23] ), .A2(\u_div/SumTmp[2][23] ), 
        .S0(quotient[2]), .Y(\u_div/PartRem[2][24] ) );
  MUX21X1_RVT U2856 ( .A1(net29741), .A2(net29939), .S0(net45600), .Y(n1072)
         );
  INVX0_RVT U2857 ( .A(\u_div/SumTmp[4][21] ), .Y(net29940) );
  INVX0_RVT U2858 ( .A(\u_div/SumTmp[6][19] ), .Y(net29942) );
  MUX21X1_RVT U2859 ( .A1(n260), .A2(n950), .S0(net46859), .Y(net29661) );
  INVX0_RVT U2860 ( .A(\u_div/SumTmp[8][17] ), .Y(net29944) );
  IBUFFX16_RVT U2861 ( .A(n1073), .Y(\u_div/PartRem[29][17] ) );
  IBUFFX16_RVT U2862 ( .A(net29976), .Y(\u_div/PartRem[28][17] ) );
  MUX21X1_RVT U2863 ( .A1(net30012), .A2(net30079), .S0(quotient[25]), .Y(
        net30033) );
  INVX0_RVT U2864 ( .A(\u_div/SumTmp[27][19] ), .Y(net30081) );
  MUX21X1_RVT U2865 ( .A1(net29956), .A2(n1081), .S0(quotient[28]), .Y(
        net29974) );
  INVX0_RVT U2866 ( .A(\u_div/SumTmp[28][18] ), .Y(n1081) );
  INVX0_RVT U2867 ( .A(\u_div/SumTmp[31][15] ), .Y(net30085) );
  INVX0_RVT U2868 ( .A(\u_div/SumTmp[33][13] ), .Y(net30087) );
  MUX21X1_RVT U2869 ( .A1(n1070), .A2(n1082), .S0(net37563), .Y(net29872) );
  MUX21X1_RVT U2870 ( .A1(n1068), .A2(n1083), .S0(net50471), .Y(n1070) );
  MUX21X1_RVT U2871 ( .A1(net44466), .A2(n1085), .S0(net37242), .Y(n1065) );
  INVX0_RVT U2872 ( .A(\u_div/SumTmp[44][2] ), .Y(net30098) );
  INVX0_RVT U2873 ( .A(\u_div/SumTmp[45][1] ), .Y(net30099) );
  NAND4X0_RVT U2874 ( .A1(n1087), .A2(n1088), .A3(n1089), .A4(n1090), .Y(n1086) );
  AND2X1_RVT U2875 ( .A1(n1091), .A2(n1092), .Y(n1090) );
  NOR3X0_RVT U2876 ( .A1(net32210), .A2(net32178), .A3(net32234), .Y(n1092) );
  NOR3X0_RVT U2877 ( .A1(b[6]), .A2(net32324), .A3(net32300), .Y(n1091) );
  AND2X1_RVT U2878 ( .A1(n1093), .A2(n1094), .Y(n1089) );
  NOR3X0_RVT U2879 ( .A1(net31814), .A2(net32352), .A3(b[2]), .Y(n1094) );
  NOR3X0_RVT U2880 ( .A1(net31896), .A2(net31844), .A3(net31872), .Y(n1093) );
  AND2X1_RVT U2881 ( .A1(n1095), .A2(n949), .Y(n1088) );
  NOR2X0_RVT U2882 ( .A1(n1096), .A2(n1097), .Y(n1087) );
  OR3X1_RVT U2883 ( .A1(net32128), .A2(net32154), .A3(n1014), .Y(n1097) );
  OR3X1_RVT U2884 ( .A1(b[14]), .A2(net32076), .A3(net32104), .Y(n1096) );
  INVX0_RVT U2885 ( .A(\u_div/SumTmp[27][18] ), .Y(net30144) );
  MUX21X1_RVT U2886 ( .A1(n1073), .A2(n1103), .S0(quotient[28]), .Y(net29975)
         );
  INVX0_RVT U2887 ( .A(\u_div/SumTmp[28][17] ), .Y(n1103) );
  MUX21X1_RVT U2888 ( .A1(net29931), .A2(net30146), .S0(net47679), .Y(n1073)
         );
  INVX0_RVT U2889 ( .A(\u_div/SumTmp[29][16] ), .Y(net30146) );
  MUX21X1_RVT U2890 ( .A1(n1071), .A2(n1104), .S0(net37563), .Y(net29873) );
  INVX0_RVT U2891 ( .A(\u_div/SumTmp[34][11] ), .Y(n1104) );
  MUX21X1_RVT U2892 ( .A1(n1069), .A2(n1105), .S0(net50471), .Y(n1071) );
  MUX21X1_RVT U2893 ( .A1(n1059), .A2(n1106), .S0(net37570), .Y(n1069) );
  INVX0_RVT U2894 ( .A(\u_div/SumTmp[36][9] ), .Y(n1106) );
  MUX21X1_RVT U2895 ( .A1(net44464), .A2(n1107), .S0(net37242), .Y(n1059) );
  INVX0_RVT U2896 ( .A(\u_div/SumTmp[37][8] ), .Y(n1107) );
  INVX0_RVT U2897 ( .A(\u_div/SumTmp[40][5] ), .Y(net30157) );
  INVX0_RVT U2898 ( .A(\u_div/SumTmp[41][4] ), .Y(net30158) );
  INVX0_RVT U2899 ( .A(\u_div/SumTmp[42][3] ), .Y(net30159) );
  INVX0_RVT U2900 ( .A(\u_div/SumTmp[44][1] ), .Y(net30161) );
  NAND4X0_RVT U2901 ( .A1(n1110), .A2(n1111), .A3(n1112), .A4(n1113), .Y(n1109) );
  NOR3X0_RVT U2902 ( .A1(net31972), .A2(net31922), .A3(net31950), .Y(n1113) );
  NOR3X0_RVT U2903 ( .A1(b[14]), .A2(net31998), .A3(net32024), .Y(n1112) );
  NOR3X0_RVT U2904 ( .A1(net32128), .A2(net32076), .A3(net32104), .Y(n1111) );
  NOR2X0_RVT U2905 ( .A1(net32154), .A2(n1114), .Y(n1110) );
  NAND4X0_RVT U2906 ( .A1(n1115), .A2(n1116), .A3(n1117), .A4(n1118), .Y(n1108) );
  NOR3X0_RVT U2907 ( .A1(net32210), .A2(net32178), .A3(net32234), .Y(n1118) );
  NOR3X0_RVT U2908 ( .A1(net32264), .A2(net32324), .A3(net32300), .Y(n1117) );
  NOR3X0_RVT U2909 ( .A1(net31814), .A2(net32352), .A3(b[2]), .Y(n1116) );
  NOR3X0_RVT U2910 ( .A1(net31896), .A2(net31844), .A3(net31872), .Y(n1115) );
  MUX21X1_RVT U2911 ( .A1(net30117), .A2(net30199), .S0(net32610), .Y(n1120)
         );
  INVX0_RVT U2912 ( .A(\u_div/SumTmp[22][22] ), .Y(net30199) );
  INVX0_RVT U2913 ( .A(\u_div/SumTmp[23][21] ), .Y(net30200) );
  MUX21X1_RVT U2914 ( .A1(n1074), .A2(n1121), .S0(quotient[28]), .Y(net29976)
         );
  INVX0_RVT U2915 ( .A(\u_div/SumTmp[28][16] ), .Y(n1121) );
  MUX21X1_RVT U2916 ( .A1(net29932), .A2(net30206), .S0(net47679), .Y(n1074)
         );
  INVX0_RVT U2917 ( .A(\u_div/SumTmp[29][15] ), .Y(net30206) );
  INVX0_RVT U2918 ( .A(\u_div/SumTmp[30][14] ), .Y(net30207) );
  INVX0_RVT U2919 ( .A(\u_div/SumTmp[31][13] ), .Y(net30208) );
  MUX21X1_RVT U2920 ( .A1(n1060), .A2(n1123), .S0(net37570), .Y(n1066) );
  INVX0_RVT U2921 ( .A(\u_div/SumTmp[36][8] ), .Y(n1123) );
  MUX21X1_RVT U2922 ( .A1(n1054), .A2(n1124), .S0(net37242), .Y(n1060) );
  INVX0_RVT U2923 ( .A(\u_div/SumTmp[37][7] ), .Y(n1124) );
  MUX21X1_RVT U2924 ( .A1(net29778), .A2(net30216), .S0(n172), .Y(net29815) );
  INVX0_RVT U2925 ( .A(\u_div/SumTmp[39][5] ), .Y(net30216) );
  INVX0_RVT U2926 ( .A(\u_div/SumTmp[40][4] ), .Y(net30217) );
  INVX0_RVT U2927 ( .A(\u_div/SumTmp[41][3] ), .Y(net30218) );
  INVX0_RVT U2928 ( .A(\u_div/SumTmp[42][2] ), .Y(net30219) );
  MUX21X1_RVT U2929 ( .A1(n1119), .A2(n1125), .S0(n192), .Y(net30245) );
  INVX0_RVT U2930 ( .A(\u_div/SumTmp[21][22] ), .Y(n1125) );
  INVX0_RVT U2931 ( .A(\u_div/SumTmp[22][21] ), .Y(net30247) );
  INVX0_RVT U2932 ( .A(\u_div/SumTmp[23][20] ), .Y(net30248) );
  INVX0_RVT U2933 ( .A(\u_div/SumTmp[27][16] ), .Y(net30252) );
  MUX21X1_RVT U2934 ( .A1(n1075), .A2(n1126), .S0(quotient[28]), .Y(net29977)
         );
  MUX21X1_RVT U2935 ( .A1(net29933), .A2(net30254), .S0(net47679), .Y(n1075)
         );
  INVX0_RVT U2936 ( .A(\u_div/SumTmp[30][13] ), .Y(net30255) );
  MUX21X1_RVT U2937 ( .A1(n1061), .A2(n1127), .S0(net37570), .Y(net29841) );
  INVX0_RVT U2938 ( .A(\u_div/SumTmp[36][7] ), .Y(n1127) );
  MUX21X1_RVT U2939 ( .A1(net29779), .A2(net30264), .S0(quotient[39]), .Y(
        net29816) );
  INVX0_RVT U2940 ( .A(\u_div/SumTmp[39][4] ), .Y(net30264) );
  INVX0_RVT U2941 ( .A(\u_div/SumTmp[40][3] ), .Y(net30265) );
  INVX0_RVT U2942 ( .A(\u_div/SumTmp[41][2] ), .Y(net30266) );
  INVX0_RVT U2943 ( .A(\u_div/SumTmp[42][1] ), .Y(net30267) );
  MUX21X1_RVT U2944 ( .A1(n951), .A2(\u_div/SumTmp[1][8] ), .S0(quotient[1]), 
        .Y(\u_div/PartRem[1][9] ) );
  INVX0_RVT U2945 ( .A(\u_div/SumTmp[6][3] ), .Y(net30289) );
  INVX0_RVT U2946 ( .A(\u_div/SumTmp[7][2] ), .Y(net30290) );
  INVX0_RVT U2947 ( .A(\u_div/SumTmp[8][1] ), .Y(net30291) );
  INVX0_RVT U2948 ( .A(\u_div/SumTmp[9][0] ), .Y(net30293) );
  MUX21X1_RVT U2949 ( .A1(\u_div/PartRem[2][7] ), .A2(\u_div/SumTmp[1][7] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][8] ) );
  MUX21X1_RVT U2950 ( .A1(n1035), .A2(n1130), .S0(n953), .Y(n1129) );
  MUX21X1_RVT U2951 ( .A1(net29730), .A2(net30296), .S0(net45582), .Y(n1035)
         );
  INVX0_RVT U2952 ( .A(\u_div/SumTmp[3][5] ), .Y(net30296) );
  INVX0_RVT U2953 ( .A(\u_div/SumTmp[5][3] ), .Y(net30298) );
  INVX0_RVT U2954 ( .A(\u_div/SumTmp[6][2] ), .Y(net30299) );
  INVX0_RVT U2955 ( .A(\u_div/SumTmp[7][1] ), .Y(net30300) );
  INVX0_RVT U2956 ( .A(\u_div/SumTmp[8][0] ), .Y(net30301) );
  MUX21X1_RVT U2957 ( .A1(\u_div/PartRem[2][6] ), .A2(\u_div/SumTmp[1][6] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][7] ) );
  MUX21X1_RVT U2958 ( .A1(n1036), .A2(n1132), .S0(quotient[2]), .Y(n1131) );
  INVX0_RVT U2959 ( .A(\u_div/SumTmp[4][3] ), .Y(net30305) );
  INVX0_RVT U2960 ( .A(\u_div/SumTmp[5][2] ), .Y(net30306) );
  INVX0_RVT U2961 ( .A(\u_div/SumTmp[6][1] ), .Y(net30307) );
  INVX0_RVT U2962 ( .A(\u_div/SumTmp[7][0] ), .Y(net30308) );
  MUX21X1_RVT U2963 ( .A1(\u_div/PartRem[2][5] ), .A2(\u_div/SumTmp[1][5] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][6] ) );
  MUX21X1_RVT U2964 ( .A1(n1037), .A2(n1134), .S0(n953), .Y(n1133) );
  MUX21X1_RVT U2965 ( .A1(net29732), .A2(net30311), .S0(net45584), .Y(n1037)
         );
  INVX0_RVT U2966 ( .A(\u_div/SumTmp[4][2] ), .Y(net30312) );
  INVX0_RVT U2967 ( .A(\u_div/SumTmp[5][1] ), .Y(net30313) );
  INVX0_RVT U2968 ( .A(\u_div/SumTmp[6][0] ), .Y(net30314) );
  MUX21X1_RVT U2969 ( .A1(\u_div/PartRem[2][4] ), .A2(\u_div/SumTmp[1][4] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][5] ) );
  MUX21X1_RVT U2970 ( .A1(n1038), .A2(n1136), .S0(n953), .Y(n1135) );
  MUX21X1_RVT U2971 ( .A1(net29733), .A2(net30317), .S0(net45601), .Y(n1038)
         );
  INVX0_RVT U2972 ( .A(\u_div/SumTmp[3][2] ), .Y(net30317) );
  INVX0_RVT U2973 ( .A(\u_div/SumTmp[4][1] ), .Y(net30318) );
  MUX21X1_RVT U2974 ( .A1(\u_div/PartRem[2][3] ), .A2(\u_div/SumTmp[1][3] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][4] ) );
  MUX21X1_RVT U2975 ( .A1(n1039), .A2(n1138), .S0(n953), .Y(n1137) );
  MUX21X1_RVT U2976 ( .A1(net29744), .A2(net30322), .S0(net45601), .Y(n1039)
         );
  INVX0_RVT U2977 ( .A(\u_div/SumTmp[3][1] ), .Y(net30322) );
  MUX21X1_RVT U2978 ( .A1(\u_div/PartRem[2][2] ), .A2(\u_div/SumTmp[1][2] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][3] ) );
  MUX21X1_RVT U2979 ( .A1(n1043), .A2(n1140), .S0(n953), .Y(n1139) );
  MUX21X1_RVT U2980 ( .A1(\u_div/PartRem[2][1] ), .A2(\u_div/SumTmp[1][1] ), 
        .S0(n1016), .Y(\u_div/PartRem[1][2] ) );
  MUX21X1_RVT U2981 ( .A1(net29742), .A2(net30331), .S0(net42514), .Y(n1041)
         );
  INVX0_RVT U2982 ( .A(\u_div/SumTmp[4][20] ), .Y(net30332) );
  INVX0_RVT U2983 ( .A(\u_div/SumTmp[6][18] ), .Y(net30334) );
  MUX21X1_RVT U2984 ( .A1(net29637), .A2(net30335), .S0(net32518), .Y(net29662) );
  INVX0_RVT U2985 ( .A(\u_div/SumTmp[7][17] ), .Y(net30335) );
  MUX21X1_RVT U2986 ( .A1(net29613), .A2(net30336), .S0(net40721), .Y(net29637) );
  INVX0_RVT U2987 ( .A(\u_div/SumTmp[8][16] ), .Y(net30336) );
  MUX21X1_RVT U2988 ( .A1(\u_div/PartRem[2][22] ), .A2(\u_div/SumTmp[1][22] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][23] ) );
  MUX21X1_RVT U2989 ( .A1(n1042), .A2(n1145), .S0(n953), .Y(n1144) );
  MUX21X1_RVT U2990 ( .A1(net29743), .A2(net30341), .S0(net45603), .Y(n1042)
         );
  INVX0_RVT U2991 ( .A(\u_div/SumTmp[3][20] ), .Y(net30341) );
  INVX0_RVT U2992 ( .A(\u_div/SumTmp[4][19] ), .Y(net30342) );
  INVX0_RVT U2993 ( .A(\u_div/SumTmp[6][17] ), .Y(net30344) );
  MUX21X1_RVT U2994 ( .A1(n1021), .A2(n1146), .S0(net46768), .Y(net29663) );
  INVX0_RVT U2995 ( .A(\u_div/SumTmp[7][16] ), .Y(n1146) );
  INVX0_RVT U2996 ( .A(\u_div/SumTmp[8][15] ), .Y(net30346) );
  MUX21X1_RVT U2997 ( .A1(\u_div/PartRem[2][21] ), .A2(\u_div/SumTmp[1][21] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][22] ) );
  MUX21X1_RVT U2998 ( .A1(net29801), .A2(n1148), .S0(n953), .Y(n1147) );
  INVX0_RVT U2999 ( .A(\u_div/SumTmp[6][16] ), .Y(net30354) );
  MUX21X1_RVT U3000 ( .A1(n1022), .A2(n1149), .S0(net32520), .Y(net29664) );
  INVX0_RVT U3001 ( .A(\u_div/SumTmp[7][15] ), .Y(n1149) );
  INVX0_RVT U3002 ( .A(\u_div/SumTmp[8][14] ), .Y(net30356) );
  MUX21X1_RVT U3003 ( .A1(\u_div/PartRem[2][20] ), .A2(\u_div/SumTmp[1][20] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][21] ) );
  MUX21X1_RVT U3004 ( .A1(n1044), .A2(n1151), .S0(n953), .Y(n1150) );
  MUX21X1_RVT U3005 ( .A1(net29746), .A2(net30361), .S0(net42523), .Y(n1044)
         );
  INVX0_RVT U3006 ( .A(\u_div/SumTmp[3][18] ), .Y(net30361) );
  INVX0_RVT U3007 ( .A(\u_div/SumTmp[4][17] ), .Y(net30362) );
  INVX0_RVT U3008 ( .A(\u_div/SumTmp[6][15] ), .Y(net30364) );
  INVX0_RVT U3009 ( .A(\u_div/SumTmp[7][14] ), .Y(n1152) );
  INVX0_RVT U3010 ( .A(\u_div/SumTmp[8][13] ), .Y(net30366) );
  MUX21X1_RVT U3011 ( .A1(\u_div/PartRem[2][19] ), .A2(\u_div/SumTmp[1][19] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][20] ) );
  MUX21X1_RVT U3012 ( .A1(n1045), .A2(n1154), .S0(n953), .Y(n1153) );
  INVX0_RVT U3013 ( .A(\u_div/SumTmp[2][18] ), .Y(n1154) );
  MUX21X1_RVT U3014 ( .A1(net29747), .A2(net30371), .S0(net45602), .Y(n1045)
         );
  INVX0_RVT U3015 ( .A(\u_div/SumTmp[3][17] ), .Y(net30371) );
  INVX0_RVT U3016 ( .A(\u_div/SumTmp[4][16] ), .Y(net30372) );
  INVX0_RVT U3017 ( .A(\u_div/SumTmp[6][14] ), .Y(net30374) );
  INVX0_RVT U3018 ( .A(\u_div/SumTmp[7][13] ), .Y(n1155) );
  INVX0_RVT U3019 ( .A(\u_div/SumTmp[8][12] ), .Y(net30376) );
  MUX21X1_RVT U3020 ( .A1(\u_div/PartRem[2][18] ), .A2(\u_div/SumTmp[1][18] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][19] ) );
  MUX21X1_RVT U3021 ( .A1(n1046), .A2(n1157), .S0(n953), .Y(n1156) );
  INVX0_RVT U3022 ( .A(\u_div/SumTmp[2][17] ), .Y(n1157) );
  MUX21X1_RVT U3023 ( .A1(net29748), .A2(net30381), .S0(net42512), .Y(n1046)
         );
  INVX0_RVT U3024 ( .A(\u_div/SumTmp[3][16] ), .Y(net30381) );
  INVX0_RVT U3025 ( .A(\u_div/SumTmp[4][15] ), .Y(net30382) );
  INVX0_RVT U3026 ( .A(\u_div/SumTmp[6][13] ), .Y(net30384) );
  INVX0_RVT U3027 ( .A(\u_div/SumTmp[7][12] ), .Y(n1158) );
  INVX0_RVT U3028 ( .A(\u_div/SumTmp[8][11] ), .Y(net30386) );
  MUX21X1_RVT U3029 ( .A1(\u_div/PartRem[2][17] ), .A2(\u_div/SumTmp[1][17] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][18] ) );
  MUX21X1_RVT U3030 ( .A1(n1047), .A2(n1160), .S0(n953), .Y(n1159) );
  INVX0_RVT U3031 ( .A(\u_div/SumTmp[2][16] ), .Y(n1160) );
  MUX21X1_RVT U3032 ( .A1(net29749), .A2(net30391), .S0(net42515), .Y(n1047)
         );
  INVX0_RVT U3033 ( .A(\u_div/SumTmp[3][15] ), .Y(net30391) );
  INVX0_RVT U3034 ( .A(\u_div/SumTmp[4][14] ), .Y(net30392) );
  INVX0_RVT U3035 ( .A(\u_div/SumTmp[6][12] ), .Y(net30394) );
  MUX21X1_RVT U3036 ( .A1(n1026), .A2(n1161), .S0(net46768), .Y(net29668) );
  INVX0_RVT U3037 ( .A(\u_div/SumTmp[7][11] ), .Y(n1161) );
  MUX21X1_RVT U3038 ( .A1(net30397), .A2(net30398), .S0(net46550), .Y(net29619) );
  MUX21X1_RVT U3039 ( .A1(\u_div/PartRem[2][16] ), .A2(\u_div/SumTmp[1][16] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][17] ) );
  MUX21X1_RVT U3040 ( .A1(n1048), .A2(n1163), .S0(n953), .Y(n1162) );
  INVX0_RVT U3041 ( .A(\u_div/SumTmp[2][15] ), .Y(n1163) );
  MUX21X1_RVT U3042 ( .A1(net29750), .A2(net30401), .S0(net42517), .Y(n1048)
         );
  INVX0_RVT U3043 ( .A(\u_div/SumTmp[3][14] ), .Y(net30401) );
  INVX0_RVT U3044 ( .A(\u_div/SumTmp[4][13] ), .Y(net30402) );
  INVX0_RVT U3045 ( .A(\u_div/SumTmp[6][11] ), .Y(net30404) );
  MUX21X1_RVT U3046 ( .A1(n1027), .A2(n1164), .S0(net46768), .Y(net29669) );
  INVX0_RVT U3047 ( .A(\u_div/SumTmp[7][10] ), .Y(n1164) );
  MUX21X1_RVT U3048 ( .A1(net29598), .A2(net30406), .S0(net40719), .Y(n1027)
         );
  INVX0_RVT U3049 ( .A(\u_div/SumTmp[8][9] ), .Y(net30406) );
  MUX21X1_RVT U3050 ( .A1(\u_div/PartRem[2][15] ), .A2(\u_div/SumTmp[1][15] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][16] ) );
  MUX21X1_RVT U3051 ( .A1(n1049), .A2(n1166), .S0(n953), .Y(n1165) );
  INVX0_RVT U3052 ( .A(\u_div/SumTmp[2][14] ), .Y(n1166) );
  MUX21X1_RVT U3053 ( .A1(net29751), .A2(net30411), .S0(net42519), .Y(n1049)
         );
  INVX0_RVT U3054 ( .A(\u_div/SumTmp[4][12] ), .Y(net30412) );
  INVX0_RVT U3055 ( .A(\u_div/SumTmp[6][10] ), .Y(net30414) );
  MUX21X1_RVT U3056 ( .A1(n1018), .A2(n1167), .S0(net46768), .Y(net29670) );
  INVX0_RVT U3057 ( .A(\u_div/SumTmp[7][9] ), .Y(n1167) );
  MUX21X1_RVT U3058 ( .A1(net29599), .A2(net30416), .S0(net40719), .Y(n1018)
         );
  INVX0_RVT U3059 ( .A(\u_div/SumTmp[8][8] ), .Y(net30416) );
  MUX21X1_RVT U3060 ( .A1(\u_div/PartRem[2][14] ), .A2(\u_div/SumTmp[1][14] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][15] ) );
  INVX0_RVT U3061 ( .A(\u_div/SumTmp[4][11] ), .Y(net30422) );
  INVX0_RVT U3062 ( .A(\u_div/SumTmp[8][7] ), .Y(net30426) );
  MUX21X1_RVT U3063 ( .A1(\u_div/PartRem[2][13] ), .A2(\u_div/SumTmp[1][13] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][14] ) );
  MUX21X1_RVT U3064 ( .A1(n1051), .A2(n1171), .S0(n953), .Y(n1170) );
  INVX0_RVT U3065 ( .A(\u_div/SumTmp[2][12] ), .Y(n1171) );
  MUX21X1_RVT U3066 ( .A1(net29753), .A2(net30431), .S0(net42520), .Y(n1051)
         );
  INVX0_RVT U3067 ( .A(\u_div/SumTmp[4][10] ), .Y(net30432) );
  INVX0_RVT U3068 ( .A(\u_div/SumTmp[5][9] ), .Y(net30433) );
  MUX21X1_RVT U3069 ( .A1(net29622), .A2(net30435), .S0(net46859), .Y(net29646) );
  INVX0_RVT U3070 ( .A(\u_div/SumTmp[7][7] ), .Y(net30435) );
  MUX21X1_RVT U3071 ( .A1(n1010), .A2(\u_div/SumTmp[1][12] ), .S0(quotient[1]), 
        .Y(\u_div/PartRem[1][13] ) );
  MUX21X1_RVT U3072 ( .A1(n995), .A2(net30441), .S0(net45588), .Y(n1052) );
  INVX0_RVT U3073 ( .A(\u_div/SumTmp[5][8] ), .Y(net30443) );
  MUX21X1_RVT U3074 ( .A1(net29623), .A2(net30445), .S0(net46859), .Y(net29647) );
  INVX0_RVT U3075 ( .A(\u_div/SumTmp[7][6] ), .Y(net30445) );
  INVX0_RVT U3076 ( .A(\u_div/SumTmp[8][5] ), .Y(net30446) );
  INVX0_RVT U3077 ( .A(\u_div/SumTmp[9][4] ), .Y(net30448) );
  MUX21X1_RVT U3078 ( .A1(n982), .A2(\u_div/SumTmp[1][11] ), .S0(quotient[1]), 
        .Y(\u_div/PartRem[1][12] ) );
  INVX0_RVT U3079 ( .A(\u_div/SumTmp[5][7] ), .Y(net30453) );
  MUX21X1_RVT U3080 ( .A1(net29624), .A2(net30455), .S0(net46859), .Y(net29648) );
  INVX0_RVT U3081 ( .A(\u_div/SumTmp[7][5] ), .Y(net30455) );
  INVX0_RVT U3082 ( .A(\u_div/SumTmp[8][4] ), .Y(net30456) );
  INVX0_RVT U3083 ( .A(\u_div/SumTmp[9][3] ), .Y(net30458) );
  INVX0_RVT U3084 ( .A(\u_div/SumTmp[2][9] ), .Y(n1173) );
  MUX21X1_RVT U3085 ( .A1(net29727), .A2(net30461), .S0(net45592), .Y(n1032)
         );
  MUX21X1_RVT U3086 ( .A1(net29649), .A2(net30464), .S0(net45257), .Y(net29674) );
  INVX0_RVT U3087 ( .A(\u_div/SumTmp[6][5] ), .Y(net30464) );
  INVX0_RVT U3088 ( .A(\u_div/SumTmp[7][4] ), .Y(net30465) );
  MUX21X1_RVT U3089 ( .A1(\u_div/PartRem[2][9] ), .A2(\u_div/SumTmp[1][9] ), 
        .S0(quotient[1]), .Y(\u_div/PartRem[1][10] ) );
  MUX21X1_RVT U3090 ( .A1(n1033), .A2(n1175), .S0(n953), .Y(n1174) );
  INVX0_RVT U3091 ( .A(\u_div/SumTmp[5][5] ), .Y(net30473) );
  INVX0_RVT U3092 ( .A(\u_div/SumTmp[6][4] ), .Y(net30474) );
  INVX0_RVT U3093 ( .A(\u_div/SumTmp[7][3] ), .Y(net30475) );
  INVX0_RVT U3094 ( .A(\u_div/SumTmp[8][2] ), .Y(net30476) );
  INVX0_RVT U3095 ( .A(\u_div/SumTmp[9][1] ), .Y(net30478) );
  MUX21X1_RVT U3096 ( .A1(net30223), .A2(net30488), .S0(net32598), .Y(net30487) );
  INVX0_RVT U3097 ( .A(\u_div/SumTmp[20][22] ), .Y(net30488) );
  INVX0_RVT U3098 ( .A(\u_div/SumTmp[21][21] ), .Y(net30489) );
  MUX21X1_RVT U3099 ( .A1(net30119), .A2(net30490), .S0(net32610), .Y(net30177) );
  INVX0_RVT U3100 ( .A(\u_div/SumTmp[22][20] ), .Y(net30490) );
  INVX0_RVT U3101 ( .A(\u_div/SumTmp[23][19] ), .Y(net30491) );
  INVX0_RVT U3102 ( .A(\u_div/SumTmp[27][15] ), .Y(net30495) );
  MUX21X1_RVT U3103 ( .A1(n1076), .A2(n1176), .S0(quotient[28]), .Y(net29978)
         );
  INVX0_RVT U3104 ( .A(\u_div/SumTmp[28][14] ), .Y(n1176) );
  MUX21X1_RVT U3105 ( .A1(net29934), .A2(net30497), .S0(net47679), .Y(n1076)
         );
  INVX0_RVT U3106 ( .A(\u_div/SumTmp[29][13] ), .Y(net30497) );
  INVX0_RVT U3107 ( .A(\u_div/SumTmp[30][12] ), .Y(net30498) );
  INVX0_RVT U3108 ( .A(\u_div/SumTmp[32][10] ), .Y(net30500) );
  MUX21X1_RVT U3109 ( .A1(n1067), .A2(n1177), .S0(net50471), .Y(net29852) );
  INVX0_RVT U3110 ( .A(\u_div/SumTmp[35][7] ), .Y(n1177) );
  MUX21X1_RVT U3111 ( .A1(n1062), .A2(n1178), .S0(net37570), .Y(n1067) );
  INVX0_RVT U3112 ( .A(\u_div/SumTmp[36][6] ), .Y(n1178) );
  MUX21X1_RVT U3113 ( .A1(n1056), .A2(n1179), .S0(net37242), .Y(n1062) );
  INVX0_RVT U3114 ( .A(\u_div/SumTmp[37][5] ), .Y(n1179) );
  INVX0_RVT U3115 ( .A(\u_div/SumTmp[38][4] ), .Y(net30506) );
  INVX0_RVT U3116 ( .A(\u_div/SumTmp[39][3] ), .Y(net30507) );
  INVX0_RVT U3117 ( .A(\u_div/SumTmp[40][2] ), .Y(net30508) );
  INVX0_RVT U3118 ( .A(\u_div/SumTmp[41][1] ), .Y(net30509) );
  MUX21X1_RVT U3119 ( .A1(net30270), .A2(net30535), .S0(net32590), .Y(net30534) );
  INVX0_RVT U3120 ( .A(\u_div/SumTmp[20][21] ), .Y(net30536) );
  INVX0_RVT U3121 ( .A(\u_div/SumTmp[21][20] ), .Y(net30537) );
  MUX21X1_RVT U3122 ( .A1(net30121), .A2(net30538), .S0(net32610), .Y(net30178) );
  INVX0_RVT U3123 ( .A(\u_div/SumTmp[22][19] ), .Y(net30538) );
  INVX0_RVT U3124 ( .A(\u_div/SumTmp[23][18] ), .Y(net30539) );
  INVX0_RVT U3125 ( .A(\u_div/SumTmp[27][14] ), .Y(net30543) );
  MUX21X1_RVT U3126 ( .A1(n1077), .A2(n1180), .S0(quotient[28]), .Y(net29979)
         );
  INVX0_RVT U3127 ( .A(\u_div/SumTmp[28][13] ), .Y(n1180) );
  MUX21X1_RVT U3128 ( .A1(net29935), .A2(net30545), .S0(net47679), .Y(n1077)
         );
  INVX0_RVT U3129 ( .A(\u_div/SumTmp[29][12] ), .Y(net30545) );
  INVX0_RVT U3130 ( .A(\u_div/SumTmp[30][11] ), .Y(net30546) );
  INVX0_RVT U3131 ( .A(\u_div/SumTmp[31][10] ), .Y(net30547) );
  INVX0_RVT U3132 ( .A(\u_div/SumTmp[32][9] ), .Y(net30548) );
  INVX0_RVT U3133 ( .A(\u_div/SumTmp[35][6] ), .Y(net30551) );
  MUX21X1_RVT U3134 ( .A1(n1063), .A2(n1181), .S0(net37570), .Y(net29843) );
  MUX21X1_RVT U3135 ( .A1(n988), .A2(n1182), .S0(net37242), .Y(n1063) );
  INVX0_RVT U3136 ( .A(\u_div/SumTmp[38][3] ), .Y(net30554) );
  INVX0_RVT U3137 ( .A(\u_div/SumTmp[39][2] ), .Y(net30555) );
  INVX0_RVT U3138 ( .A(\u_div/SumTmp[40][1] ), .Y(net30556) );
  MUX21X1_RVT U3139 ( .A1(net30271), .A2(net30583), .S0(net32590), .Y(net30512) );
  INVX0_RVT U3140 ( .A(\u_div/SumTmp[20][20] ), .Y(net30584) );
  INVX0_RVT U3141 ( .A(\u_div/SumTmp[21][19] ), .Y(net30585) );
  MUX21X1_RVT U3142 ( .A1(net30122), .A2(net30586), .S0(net32610), .Y(net30180) );
  INVX0_RVT U3143 ( .A(\u_div/SumTmp[22][18] ), .Y(net30586) );
  INVX0_RVT U3144 ( .A(\u_div/SumTmp[23][17] ), .Y(net30587) );
  INVX0_RVT U3145 ( .A(\u_div/SumTmp[27][13] ), .Y(net30591) );
  MUX21X1_RVT U3146 ( .A1(n1078), .A2(n1183), .S0(quotient[28]), .Y(net29980)
         );
  MUX21X1_RVT U3147 ( .A1(net29936), .A2(net30593), .S0(net47679), .Y(n1078)
         );
  INVX0_RVT U3148 ( .A(\u_div/SumTmp[29][11] ), .Y(net30593) );
  INVX0_RVT U3149 ( .A(\u_div/SumTmp[30][10] ), .Y(net30594) );
  INVX0_RVT U3150 ( .A(\u_div/SumTmp[31][9] ), .Y(net30595) );
  INVX0_RVT U3151 ( .A(\u_div/SumTmp[32][8] ), .Y(net30596) );
  INVX0_RVT U3152 ( .A(\u_div/SumTmp[33][7] ), .Y(net30597) );
  MUX21X1_RVT U3153 ( .A1(n1064), .A2(n1184), .S0(net37570), .Y(net29844) );
  INVX0_RVT U3154 ( .A(\u_div/SumTmp[36][4] ), .Y(n1184) );
  MUX21X1_RVT U3155 ( .A1(n1058), .A2(n1185), .S0(net37242), .Y(n1064) );
  INVX0_RVT U3156 ( .A(\u_div/SumTmp[37][3] ), .Y(n1185) );
  MUX21X1_RVT U3157 ( .A1(net29782), .A2(net30603), .S0(n172), .Y(net29819) );
  INVX0_RVT U3158 ( .A(\u_div/SumTmp[39][1] ), .Y(net30603) );
  MUX21X1_RVT U3159 ( .A1(net30559), .A2(net30629), .S0(n158), .Y(net30628) );
  INVX0_RVT U3160 ( .A(\u_div/SumTmp[20][19] ), .Y(net30632) );
  INVX0_RVT U3161 ( .A(\u_div/SumTmp[21][18] ), .Y(net30633) );
  INVX0_RVT U3162 ( .A(\u_div/SumTmp[22][17] ), .Y(net30634) );
  INVX0_RVT U3163 ( .A(\u_div/SumTmp[23][16] ), .Y(net30635) );
  MUX21X1_RVT U3164 ( .A1(n1079), .A2(n1186), .S0(quotient[28]), .Y(net29981)
         );
  MUX21X1_RVT U3165 ( .A1(net29937), .A2(net30641), .S0(net47679), .Y(n1079)
         );
  INVX0_RVT U3166 ( .A(\u_div/SumTmp[29][10] ), .Y(net30641) );
  INVX0_RVT U3167 ( .A(\u_div/SumTmp[30][9] ), .Y(net30642) );
  INVX0_RVT U3168 ( .A(\u_div/SumTmp[31][8] ), .Y(net30643) );
  INVX0_RVT U3169 ( .A(\u_div/SumTmp[32][7] ), .Y(net30644) );
  INVX0_RVT U3170 ( .A(\u_div/SumTmp[33][6] ), .Y(net30645) );
  MUX21X1_RVT U3171 ( .A1(net30606), .A2(net30676), .S0(n17), .Y(net30675) );
  INVX0_RVT U3172 ( .A(\u_div/SumTmp[16][22] ), .Y(net30676) );
  INVX0_RVT U3173 ( .A(\u_div/SumTmp[20][18] ), .Y(net30680) );
  INVX0_RVT U3174 ( .A(\u_div/SumTmp[21][17] ), .Y(net30681) );
  MUX21X1_RVT U3175 ( .A1(net30124), .A2(n1187), .S0(net32610), .Y(net30182)
         );
  INVX0_RVT U3176 ( .A(\u_div/SumTmp[22][16] ), .Y(n1187) );
  MUX21X1_RVT U3177 ( .A1(net30063), .A2(net30683), .S0(quotient[23]), .Y(
        net30124) );
  INVX0_RVT U3178 ( .A(\u_div/SumTmp[23][15] ), .Y(net30683) );
  MUX21X1_RVT U3179 ( .A1(n1080), .A2(n1188), .S0(quotient[28]), .Y(net29982)
         );
  INVX0_RVT U3180 ( .A(\u_div/SumTmp[28][10] ), .Y(n1188) );
  MUX21X1_RVT U3181 ( .A1(net29921), .A2(net30689), .S0(net47679), .Y(n1080)
         );
  INVX0_RVT U3182 ( .A(\u_div/SumTmp[29][9] ), .Y(net30689) );
  INVX0_RVT U3183 ( .A(\u_div/SumTmp[30][8] ), .Y(net30690) );
  INVX0_RVT U3184 ( .A(\u_div/SumTmp[31][7] ), .Y(net30691) );
  INVX0_RVT U3185 ( .A(\u_div/SumTmp[32][6] ), .Y(net30692) );
  INVX0_RVT U3186 ( .A(\u_div/SumTmp[33][5] ), .Y(net30693) );
  INVX0_RVT U3187 ( .A(\u_div/SumTmp[34][4] ), .Y(net30694) );
  INVX0_RVT U3188 ( .A(\u_div/SumTmp[35][3] ), .Y(net30695) );
  INVX0_RVT U3189 ( .A(\u_div/SumTmp[36][2] ), .Y(net30696) );
  MUX21X1_RVT U3190 ( .A1(\u_div/PartRem[15][23] ), .A2(\u_div/SumTmp[14][23] ), .S0(net32560), .Y(\u_div/PartRem[14][24] ) );
  MUX21X1_RVT U3191 ( .A1(net30653), .A2(net30723), .S0(n56), .Y(n1191) );
  INVX0_RVT U3192 ( .A(\u_div/SumTmp[16][21] ), .Y(net30724) );
  INVX0_RVT U3193 ( .A(\u_div/SumTmp[20][17] ), .Y(net30728) );
  INVX0_RVT U3194 ( .A(\u_div/SumTmp[21][16] ), .Y(net30729) );
  MUX21X1_RVT U3195 ( .A1(n1098), .A2(n1192), .S0(net32610), .Y(net30183) );
  INVX0_RVT U3196 ( .A(\u_div/SumTmp[22][15] ), .Y(n1192) );
  MUX21X1_RVT U3197 ( .A1(net30064), .A2(net30731), .S0(quotient[23]), .Y(
        n1098) );
  INVX0_RVT U3198 ( .A(\u_div/SumTmp[23][14] ), .Y(net30731) );
  INVX0_RVT U3199 ( .A(\u_div/SumTmp[24][13] ), .Y(net30732) );
  INVX0_RVT U3200 ( .A(\u_div/SumTmp[29][8] ), .Y(net30737) );
  INVX0_RVT U3201 ( .A(\u_div/SumTmp[30][7] ), .Y(net30738) );
  INVX0_RVT U3202 ( .A(\u_div/SumTmp[31][6] ), .Y(net30739) );
  INVX0_RVT U3203 ( .A(\u_div/SumTmp[32][5] ), .Y(net30740) );
  INVX0_RVT U3204 ( .A(\u_div/SumTmp[33][4] ), .Y(net30741) );
  INVX0_RVT U3205 ( .A(\u_div/SumTmp[34][3] ), .Y(net30742) );
  INVX0_RVT U3206 ( .A(\u_div/SumTmp[35][2] ), .Y(net30743) );
  INVX0_RVT U3207 ( .A(\u_div/SumTmp[36][1] ), .Y(net30744) );
  MUX21X1_RVT U3208 ( .A1(\u_div/PartRem[14][23] ), .A2(\u_div/SumTmp[13][23] ), .S0(net42408), .Y(\u_div/PartRem[13][24] ) );
  MUX21X1_RVT U3209 ( .A1(n1189), .A2(n1195), .S0(net32560), .Y(n1194) );
  MUX21X1_RVT U3210 ( .A1(net30654), .A2(net30771), .S0(quotient[15]), .Y(
        n1189) );
  INVX0_RVT U3211 ( .A(\u_div/SumTmp[16][20] ), .Y(net30772) );
  INVX0_RVT U3212 ( .A(\u_div/SumTmp[17][19] ), .Y(net30773) );
  INVX0_RVT U3213 ( .A(\u_div/SumTmp[21][15] ), .Y(net30777) );
  MUX21X1_RVT U3214 ( .A1(n1099), .A2(n1196), .S0(net32610), .Y(net30184) );
  INVX0_RVT U3215 ( .A(\u_div/SumTmp[22][14] ), .Y(n1196) );
  MUX21X1_RVT U3216 ( .A1(net30065), .A2(net30779), .S0(quotient[23]), .Y(
        n1099) );
  INVX0_RVT U3217 ( .A(\u_div/SumTmp[23][13] ), .Y(net30779) );
  INVX0_RVT U3218 ( .A(\u_div/SumTmp[24][12] ), .Y(net30780) );
  INVX0_RVT U3219 ( .A(\u_div/SumTmp[26][10] ), .Y(net30782) );
  INVX0_RVT U3220 ( .A(\u_div/SumTmp[29][7] ), .Y(net30785) );
  INVX0_RVT U3221 ( .A(\u_div/SumTmp[30][6] ), .Y(net30786) );
  INVX0_RVT U3222 ( .A(\u_div/SumTmp[32][4] ), .Y(net30788) );
  INVX0_RVT U3223 ( .A(\u_div/SumTmp[33][3] ), .Y(net30789) );
  INVX0_RVT U3224 ( .A(\u_div/SumTmp[34][2] ), .Y(net30790) );
  INVX0_RVT U3225 ( .A(\u_div/SumTmp[35][1] ), .Y(net30791) );
  MUX21X1_RVT U3226 ( .A1(n1190), .A2(n1198), .S0(net32560), .Y(n1193) );
  INVX0_RVT U3227 ( .A(\u_div/SumTmp[14][21] ), .Y(n1198) );
  MUX21X1_RVT U3228 ( .A1(net30655), .A2(net30819), .S0(n52), .Y(n1190) );
  INVX0_RVT U3229 ( .A(\u_div/SumTmp[16][19] ), .Y(net30820) );
  INVX0_RVT U3230 ( .A(\u_div/SumTmp[21][14] ), .Y(net30825) );
  MUX21X1_RVT U3231 ( .A1(n1100), .A2(n1199), .S0(net32608), .Y(net30185) );
  INVX0_RVT U3232 ( .A(\u_div/SumTmp[22][13] ), .Y(n1199) );
  MUX21X1_RVT U3233 ( .A1(net30066), .A2(net30827), .S0(quotient[23]), .Y(
        n1100) );
  INVX0_RVT U3234 ( .A(\u_div/SumTmp[23][12] ), .Y(net30827) );
  INVX0_RVT U3235 ( .A(\u_div/SumTmp[24][11] ), .Y(net30828) );
  INVX0_RVT U3236 ( .A(\u_div/SumTmp[27][8] ), .Y(net30831) );
  INVX0_RVT U3237 ( .A(\u_div/SumTmp[29][6] ), .Y(net30833) );
  INVX0_RVT U3238 ( .A(\u_div/SumTmp[30][5] ), .Y(net30834) );
  INVX0_RVT U3239 ( .A(\u_div/SumTmp[31][4] ), .Y(net30835) );
  INVX0_RVT U3240 ( .A(\u_div/SumTmp[32][3] ), .Y(net30836) );
  INVX0_RVT U3241 ( .A(\u_div/SumTmp[33][2] ), .Y(net30837) );
  INVX0_RVT U3242 ( .A(\u_div/SumTmp[34][1] ), .Y(net30838) );
  MUX21X1_RVT U3243 ( .A1(net30794), .A2(net30864), .S0(net32548), .Y(net30863) );
  INVX0_RVT U3244 ( .A(\u_div/SumTmp[13][21] ), .Y(net30865) );
  MUX21X1_RVT U3245 ( .A1(net30702), .A2(net30866), .S0(net32560), .Y(net30748) );
  INVX0_RVT U3246 ( .A(\u_div/SumTmp[14][20] ), .Y(net30866) );
  MUX21X1_RVT U3247 ( .A1(net30657), .A2(net30867), .S0(n50), .Y(net30702) );
  INVX0_RVT U3248 ( .A(\u_div/SumTmp[16][18] ), .Y(net30868) );
  INVX0_RVT U3249 ( .A(\u_div/SumTmp[18][16] ), .Y(net30870) );
  INVX0_RVT U3250 ( .A(\u_div/SumTmp[19][15] ), .Y(net30871) );
  INVX0_RVT U3251 ( .A(\u_div/SumTmp[21][13] ), .Y(net30873) );
  MUX21X1_RVT U3252 ( .A1(n1101), .A2(n1200), .S0(net32608), .Y(net30186) );
  INVX0_RVT U3253 ( .A(\u_div/SumTmp[22][12] ), .Y(n1200) );
  MUX21X1_RVT U3254 ( .A1(net30067), .A2(net30875), .S0(quotient[23]), .Y(
        n1101) );
  INVX0_RVT U3255 ( .A(\u_div/SumTmp[23][11] ), .Y(net30875) );
  INVX0_RVT U3256 ( .A(\u_div/SumTmp[24][10] ), .Y(net30876) );
  INVX0_RVT U3257 ( .A(\u_div/SumTmp[27][7] ), .Y(net30879) );
  INVX0_RVT U3258 ( .A(\u_div/SumTmp[29][5] ), .Y(net30881) );
  INVX0_RVT U3259 ( .A(\u_div/SumTmp[30][4] ), .Y(net30882) );
  INVX0_RVT U3260 ( .A(\u_div/SumTmp[31][3] ), .Y(net30883) );
  INVX0_RVT U3261 ( .A(\u_div/SumTmp[32][2] ), .Y(net30884) );
  INVX0_RVT U3262 ( .A(\u_div/SumTmp[33][1] ), .Y(net30885) );
  INVX0_RVT U3263 ( .A(\u_div/SumTmp[10][8] ), .Y(net30902) );
  INVX0_RVT U3264 ( .A(\u_div/SumTmp[11][7] ), .Y(net30903) );
  INVX0_RVT U3265 ( .A(\u_div/SumTmp[12][6] ), .Y(net30904) );
  INVX0_RVT U3266 ( .A(\u_div/SumTmp[13][5] ), .Y(net30905) );
  INVX0_RVT U3267 ( .A(\u_div/SumTmp[14][4] ), .Y(net30906) );
  INVX0_RVT U3268 ( .A(\u_div/SumTmp[15][3] ), .Y(net30907) );
  INVX0_RVT U3269 ( .A(\u_div/SumTmp[17][1] ), .Y(net30909) );
  INVX0_RVT U3270 ( .A(\u_div/SumTmp[18][0] ), .Y(net30910) );
  INVX0_RVT U3271 ( .A(\u_div/SumTmp[10][7] ), .Y(net30911) );
  INVX0_RVT U3272 ( .A(\u_div/SumTmp[11][6] ), .Y(net30912) );
  INVX0_RVT U3273 ( .A(\u_div/SumTmp[12][5] ), .Y(net30913) );
  INVX0_RVT U3274 ( .A(\u_div/SumTmp[13][4] ), .Y(net30914) );
  INVX0_RVT U3275 ( .A(\u_div/SumTmp[15][2] ), .Y(net30916) );
  INVX0_RVT U3276 ( .A(\u_div/SumTmp[10][6] ), .Y(net30919) );
  INVX0_RVT U3277 ( .A(\u_div/SumTmp[11][5] ), .Y(net30920) );
  INVX0_RVT U3278 ( .A(\u_div/SumTmp[12][4] ), .Y(net30921) );
  INVX0_RVT U3279 ( .A(\u_div/SumTmp[13][3] ), .Y(net30922) );
  INVX0_RVT U3280 ( .A(\u_div/SumTmp[14][2] ), .Y(net30923) );
  INVX0_RVT U3281 ( .A(\u_div/SumTmp[15][1] ), .Y(net30924) );
  INVX0_RVT U3282 ( .A(\u_div/SumTmp[16][0] ), .Y(net30925) );
  INVX0_RVT U3283 ( .A(\u_div/SumTmp[10][5] ), .Y(net30926) );
  INVX0_RVT U3284 ( .A(\u_div/SumTmp[11][4] ), .Y(net30927) );
  INVX0_RVT U3285 ( .A(\u_div/SumTmp[12][3] ), .Y(net30928) );
  INVX0_RVT U3286 ( .A(\u_div/SumTmp[13][2] ), .Y(net30929) );
  INVX0_RVT U3287 ( .A(\u_div/SumTmp[14][1] ), .Y(net30930) );
  INVX0_RVT U3288 ( .A(\u_div/SumTmp[15][0] ), .Y(net30931) );
  INVX0_RVT U3289 ( .A(\u_div/SumTmp[11][3] ), .Y(net30933) );
  INVX0_RVT U3290 ( .A(\u_div/SumTmp[12][2] ), .Y(net30934) );
  INVX0_RVT U3291 ( .A(\u_div/SumTmp[13][1] ), .Y(net30935) );
  INVX0_RVT U3292 ( .A(\u_div/SumTmp[14][0] ), .Y(net30936) );
  INVX0_RVT U3293 ( .A(\u_div/SumTmp[10][3] ), .Y(net30937) );
  INVX0_RVT U3294 ( .A(\u_div/SumTmp[11][2] ), .Y(net30938) );
  INVX0_RVT U3295 ( .A(\u_div/SumTmp[12][1] ), .Y(net30939) );
  INVX0_RVT U3296 ( .A(\u_div/SumTmp[13][0] ), .Y(net30940) );
  INVX0_RVT U3297 ( .A(\u_div/SumTmp[10][2] ), .Y(net30941) );
  INVX0_RVT U3298 ( .A(\u_div/SumTmp[11][1] ), .Y(net30942) );
  INVX0_RVT U3299 ( .A(\u_div/SumTmp[12][0] ), .Y(net30943) );
  INVX0_RVT U3300 ( .A(\u_div/SumTmp[10][1] ), .Y(net30944) );
  INVX0_RVT U3301 ( .A(\u_div/SumTmp[11][0] ), .Y(net30945) );
  INVX0_RVT U3302 ( .A(\u_div/SumTmp[16][17] ), .Y(net30952) );
  INVX0_RVT U3303 ( .A(\u_div/SumTmp[17][16] ), .Y(net30953) );
  INVX0_RVT U3304 ( .A(\u_div/SumTmp[18][15] ), .Y(net30954) );
  INVX0_RVT U3305 ( .A(\u_div/SumTmp[19][14] ), .Y(net30955) );
  INVX0_RVT U3306 ( .A(\u_div/SumTmp[21][12] ), .Y(net30957) );
  MUX21X1_RVT U3307 ( .A1(n1102), .A2(n1201), .S0(net32608), .Y(net30187) );
  INVX0_RVT U3308 ( .A(\u_div/SumTmp[22][11] ), .Y(n1201) );
  INVX0_RVT U3309 ( .A(\u_div/SumTmp[23][10] ), .Y(net30959) );
  INVX0_RVT U3310 ( .A(\u_div/SumTmp[25][8] ), .Y(net30961) );
  INVX0_RVT U3311 ( .A(\u_div/SumTmp[27][6] ), .Y(net30963) );
  INVX0_RVT U3312 ( .A(\u_div/SumTmp[29][4] ), .Y(net30965) );
  INVX0_RVT U3313 ( .A(\u_div/SumTmp[30][3] ), .Y(net30966) );
  INVX0_RVT U3314 ( .A(\u_div/SumTmp[31][2] ), .Y(net30967) );
  INVX0_RVT U3315 ( .A(\u_div/SumTmp[32][1] ), .Y(net30968) );
  MUX21X1_RVT U3316 ( .A1(net30888), .A2(net30972), .S0(net32538), .Y(n1202)
         );
  INVX0_RVT U3317 ( .A(\u_div/SumTmp[11][21] ), .Y(net30973) );
  INVX0_RVT U3318 ( .A(\u_div/SumTmp[13][19] ), .Y(net30975) );
  MUX21X1_RVT U3319 ( .A1(net30613), .A2(net30978), .S0(n19), .Y(net30659) );
  INVX0_RVT U3320 ( .A(\u_div/SumTmp[17][15] ), .Y(net30979) );
  INVX0_RVT U3321 ( .A(\u_div/SumTmp[18][14] ), .Y(net30980) );
  INVX0_RVT U3322 ( .A(\u_div/SumTmp[19][13] ), .Y(net30981) );
  INVX0_RVT U3323 ( .A(\u_div/SumTmp[22][10] ), .Y(net30984) );
  MUX21X1_RVT U3324 ( .A1(net30047), .A2(net30985), .S0(quotient[23]), .Y(
        net30130) );
  INVX0_RVT U3325 ( .A(\u_div/SumTmp[23][9] ), .Y(net30985) );
  INVX0_RVT U3326 ( .A(\u_div/SumTmp[25][7] ), .Y(net30987) );
  INVX0_RVT U3327 ( .A(\u_div/SumTmp[26][6] ), .Y(net30988) );
  INVX0_RVT U3328 ( .A(\u_div/SumTmp[27][5] ), .Y(net30989) );
  INVX0_RVT U3329 ( .A(\u_div/SumTmp[29][3] ), .Y(net30991) );
  INVX0_RVT U3330 ( .A(\u_div/SumTmp[31][1] ), .Y(net30993) );
  MUX21X1_RVT U3331 ( .A1(net30889), .A2(net30996), .S0(net32536), .Y(n1019)
         );
  INVX0_RVT U3332 ( .A(\u_div/SumTmp[11][20] ), .Y(net30997) );
  INVX0_RVT U3333 ( .A(\u_div/SumTmp[13][18] ), .Y(net30999) );
  INVX0_RVT U3334 ( .A(\u_div/SumTmp[16][15] ), .Y(net31002) );
  INVX0_RVT U3335 ( .A(\u_div/SumTmp[17][14] ), .Y(net31003) );
  INVX0_RVT U3336 ( .A(\u_div/SumTmp[18][13] ), .Y(net31004) );
  INVX0_RVT U3337 ( .A(\u_div/SumTmp[19][12] ), .Y(net31005) );
  INVX0_RVT U3338 ( .A(\u_div/SumTmp[20][11] ), .Y(net31006) );
  INVX0_RVT U3339 ( .A(\u_div/SumTmp[22][9] ), .Y(net31008) );
  MUX21X1_RVT U3340 ( .A1(net30048), .A2(net31009), .S0(quotient[23]), .Y(
        net30069) );
  INVX0_RVT U3341 ( .A(\u_div/SumTmp[23][8] ), .Y(net31009) );
  INVX0_RVT U3342 ( .A(\u_div/SumTmp[24][7] ), .Y(net31010) );
  INVX0_RVT U3343 ( .A(\u_div/SumTmp[27][4] ), .Y(net31013) );
  INVX0_RVT U3344 ( .A(\u_div/SumTmp[29][2] ), .Y(net31015) );
  MUX21X1_RVT U3345 ( .A1(net30890), .A2(net31019), .S0(net32538), .Y(net29655) );
  INVX0_RVT U3346 ( .A(\u_div/SumTmp[11][19] ), .Y(net31020) );
  INVX0_RVT U3347 ( .A(\u_div/SumTmp[17][13] ), .Y(net31026) );
  INVX0_RVT U3348 ( .A(\u_div/SumTmp[18][12] ), .Y(net31027) );
  INVX0_RVT U3349 ( .A(\u_div/SumTmp[19][11] ), .Y(net31028) );
  INVX0_RVT U3350 ( .A(\u_div/SumTmp[20][10] ), .Y(net31029) );
  INVX0_RVT U3351 ( .A(\u_div/SumTmp[22][8] ), .Y(net31031) );
  MUX21X1_RVT U3352 ( .A1(net30049), .A2(net31032), .S0(quotient[23]), .Y(
        net30070) );
  INVX0_RVT U3353 ( .A(\u_div/SumTmp[23][7] ), .Y(net31032) );
  INVX0_RVT U3354 ( .A(\u_div/SumTmp[24][6] ), .Y(net31033) );
  INVX0_RVT U3355 ( .A(\u_div/SumTmp[25][5] ), .Y(net31034) );
  INVX0_RVT U3356 ( .A(\u_div/SumTmp[26][4] ), .Y(net31035) );
  INVX0_RVT U3357 ( .A(\u_div/SumTmp[29][1] ), .Y(net31038) );
  MUX21X1_RVT U3358 ( .A1(net30892), .A2(net31041), .S0(net32538), .Y(net29682) );
  INVX0_RVT U3359 ( .A(\u_div/SumTmp[12][17] ), .Y(net31043) );
  INVX0_RVT U3360 ( .A(\u_div/SumTmp[13][16] ), .Y(net31044) );
  INVX0_RVT U3361 ( .A(\u_div/SumTmp[17][12] ), .Y(net31048) );
  INVX0_RVT U3362 ( .A(\u_div/SumTmp[18][11] ), .Y(net31049) );
  INVX0_RVT U3363 ( .A(\u_div/SumTmp[19][10] ), .Y(net31050) );
  INVX0_RVT U3364 ( .A(\u_div/SumTmp[20][9] ), .Y(net31051) );
  INVX0_RVT U3365 ( .A(\u_div/SumTmp[22][7] ), .Y(net31053) );
  MUX21X1_RVT U3366 ( .A1(net30050), .A2(net31054), .S0(quotient[23]), .Y(
        net30071) );
  INVX0_RVT U3367 ( .A(\u_div/SumTmp[23][6] ), .Y(net31054) );
  INVX0_RVT U3368 ( .A(\u_div/SumTmp[24][5] ), .Y(net31055) );
  INVX0_RVT U3369 ( .A(\u_div/SumTmp[27][2] ), .Y(net31058) );
  MUX21X1_RVT U3370 ( .A1(net30893), .A2(net31063), .S0(net32538), .Y(net29710) );
  INVX0_RVT U3371 ( .A(\u_div/SumTmp[11][17] ), .Y(net31064) );
  INVX0_RVT U3372 ( .A(\u_div/SumTmp[15][13] ), .Y(net31068) );
  INVX0_RVT U3373 ( .A(\u_div/SumTmp[17][11] ), .Y(net31070) );
  INVX0_RVT U3374 ( .A(\u_div/SumTmp[18][10] ), .Y(net31071) );
  INVX0_RVT U3375 ( .A(\u_div/SumTmp[19][9] ), .Y(net31072) );
  INVX0_RVT U3376 ( .A(\u_div/SumTmp[20][8] ), .Y(net31073) );
  INVX0_RVT U3377 ( .A(\u_div/SumTmp[22][6] ), .Y(net31075) );
  MUX21X1_RVT U3378 ( .A1(net30051), .A2(net31076), .S0(quotient[23]), .Y(
        net30072) );
  INVX0_RVT U3379 ( .A(\u_div/SumTmp[23][5] ), .Y(net31076) );
  INVX0_RVT U3380 ( .A(\u_div/SumTmp[25][3] ), .Y(net31078) );
  INVX0_RVT U3381 ( .A(\u_div/SumTmp[26][2] ), .Y(net31079) );
  INVX0_RVT U3382 ( .A(\u_div/SumTmp[27][1] ), .Y(net31080) );
  INVX0_RVT U3383 ( .A(\u_div/SumTmp[11][16] ), .Y(net31084) );
  INVX0_RVT U3384 ( .A(\u_div/SumTmp[13][14] ), .Y(net31086) );
  INVX0_RVT U3385 ( .A(\u_div/SumTmp[15][12] ), .Y(net31088) );
  INVX0_RVT U3386 ( .A(\u_div/SumTmp[17][10] ), .Y(net31090) );
  INVX0_RVT U3387 ( .A(\u_div/SumTmp[18][9] ), .Y(net31091) );
  INVX0_RVT U3388 ( .A(\u_div/SumTmp[19][8] ), .Y(net31092) );
  INVX0_RVT U3389 ( .A(\u_div/SumTmp[20][7] ), .Y(net31093) );
  INVX0_RVT U3390 ( .A(\u_div/SumTmp[23][4] ), .Y(net31096) );
  INVX0_RVT U3391 ( .A(\u_div/SumTmp[25][2] ), .Y(net31098) );
  INVX0_RVT U3392 ( .A(\u_div/SumTmp[26][1] ), .Y(net31099) );
  INVX0_RVT U3393 ( .A(\u_div/SumTmp[11][15] ), .Y(net31103) );
  INVX0_RVT U3394 ( .A(\u_div/SumTmp[17][9] ), .Y(net31109) );
  INVX0_RVT U3395 ( .A(\u_div/SumTmp[18][8] ), .Y(net31110) );
  INVX0_RVT U3396 ( .A(\u_div/SumTmp[19][7] ), .Y(net31111) );
  INVX0_RVT U3397 ( .A(\u_div/SumTmp[20][6] ), .Y(net31112) );
  INVX0_RVT U3398 ( .A(\u_div/SumTmp[21][5] ), .Y(net31113) );
  INVX0_RVT U3399 ( .A(\u_div/SumTmp[23][3] ), .Y(net31115) );
  INVX0_RVT U3400 ( .A(\u_div/SumTmp[25][1] ), .Y(net31117) );
  INVX0_RVT U3401 ( .A(\u_div/SumTmp[12][13] ), .Y(net31122) );
  INVX0_RVT U3402 ( .A(\u_div/SumTmp[15][10] ), .Y(net31125) );
  INVX0_RVT U3403 ( .A(\u_div/SumTmp[17][8] ), .Y(net31127) );
  INVX0_RVT U3404 ( .A(\u_div/SumTmp[18][7] ), .Y(net31128) );
  INVX0_RVT U3405 ( .A(\u_div/SumTmp[19][6] ), .Y(net31129) );
  INVX0_RVT U3406 ( .A(\u_div/SumTmp[20][5] ), .Y(net31130) );
  INVX0_RVT U3407 ( .A(\u_div/SumTmp[21][4] ), .Y(net31131) );
  INVX0_RVT U3408 ( .A(\u_div/SumTmp[22][3] ), .Y(net31132) );
  INVX0_RVT U3409 ( .A(\u_div/SumTmp[23][2] ), .Y(net31133) );
  INVX0_RVT U3410 ( .A(\u_div/SumTmp[11][13] ), .Y(net31138) );
  INVX0_RVT U3411 ( .A(\u_div/SumTmp[12][12] ), .Y(net31139) );
  INVX0_RVT U3412 ( .A(\u_div/SumTmp[14][10] ), .Y(net31141) );
  INVX0_RVT U3413 ( .A(\u_div/SumTmp[15][9] ), .Y(net31142) );
  INVX0_RVT U3414 ( .A(\u_div/SumTmp[17][7] ), .Y(net31144) );
  INVX0_RVT U3415 ( .A(\u_div/SumTmp[18][6] ), .Y(net31145) );
  INVX0_RVT U3416 ( .A(\u_div/SumTmp[19][5] ), .Y(net31146) );
  INVX0_RVT U3417 ( .A(\u_div/SumTmp[20][4] ), .Y(net31147) );
  INVX0_RVT U3418 ( .A(\u_div/SumTmp[21][3] ), .Y(net31148) );
  INVX0_RVT U3419 ( .A(\u_div/SumTmp[22][2] ), .Y(net31149) );
  INVX0_RVT U3420 ( .A(\u_div/SumTmp[23][1] ), .Y(net31150) );
  INVX0_RVT U3421 ( .A(\u_div/SumTmp[11][12] ), .Y(net31154) );
  INVX0_RVT U3422 ( .A(\u_div/SumTmp[15][8] ), .Y(net31158) );
  INVX0_RVT U3423 ( .A(\u_div/SumTmp[17][6] ), .Y(net31160) );
  INVX0_RVT U3424 ( .A(\u_div/SumTmp[18][5] ), .Y(net31161) );
  INVX0_RVT U3425 ( .A(\u_div/SumTmp[19][4] ), .Y(net31162) );
  INVX0_RVT U3426 ( .A(\u_div/SumTmp[20][3] ), .Y(net31163) );
  INVX0_RVT U3427 ( .A(\u_div/SumTmp[21][2] ), .Y(net31164) );
  INVX0_RVT U3428 ( .A(\u_div/SumTmp[22][1] ), .Y(net31165) );
  MUX21X1_RVT U3429 ( .A1(net30807), .A2(net31170), .S0(quotient[12]), .Y(
        net30853) );
  INVX0_RVT U3430 ( .A(\u_div/SumTmp[12][10] ), .Y(net31170) );
  INVX0_RVT U3431 ( .A(\u_div/SumTmp[17][5] ), .Y(net31175) );
  INVX0_RVT U3432 ( .A(\u_div/SumTmp[18][4] ), .Y(net31176) );
  INVX0_RVT U3433 ( .A(\u_div/SumTmp[19][3] ), .Y(net31177) );
  INVX0_RVT U3434 ( .A(\u_div/SumTmp[20][2] ), .Y(net31178) );
  INVX0_RVT U3435 ( .A(\u_div/SumTmp[21][1] ), .Y(net31179) );
  INVX0_RVT U3436 ( .A(\u_div/SumTmp[22][0] ), .Y(net31180) );
  INVX0_RVT U3437 ( .A(\u_div/SumTmp[10][11] ), .Y(net31181) );
  INVX0_RVT U3438 ( .A(\u_div/SumTmp[11][10] ), .Y(net31182) );
  INVX0_RVT U3439 ( .A(\u_div/SumTmp[12][9] ), .Y(net31183) );
  INVX0_RVT U3440 ( .A(\u_div/SumTmp[14][7] ), .Y(net31185) );
  INVX0_RVT U3441 ( .A(\u_div/SumTmp[15][6] ), .Y(net31186) );
  INVX0_RVT U3442 ( .A(\u_div/SumTmp[17][4] ), .Y(net31188) );
  INVX0_RVT U3443 ( .A(\u_div/SumTmp[18][3] ), .Y(net31189) );
  INVX0_RVT U3444 ( .A(\u_div/SumTmp[19][2] ), .Y(net31190) );
  INVX0_RVT U3445 ( .A(\u_div/SumTmp[20][1] ), .Y(net31191) );
  INVX0_RVT U3446 ( .A(\u_div/SumTmp[21][0] ), .Y(net31192) );
  INVX0_RVT U3447 ( .A(\u_div/SumTmp[10][10] ), .Y(net31193) );
  INVX0_RVT U3448 ( .A(\u_div/SumTmp[11][9] ), .Y(net31194) );
  INVX0_RVT U3449 ( .A(\u_div/SumTmp[12][8] ), .Y(net31195) );
  INVX0_RVT U3450 ( .A(\u_div/SumTmp[15][5] ), .Y(net31198) );
  INVX0_RVT U3451 ( .A(\u_div/SumTmp[17][3] ), .Y(net31200) );
  INVX0_RVT U3452 ( .A(\u_div/SumTmp[18][2] ), .Y(net31201) );
  INVX0_RVT U3453 ( .A(\u_div/SumTmp[19][1] ), .Y(net31202) );
  INVX0_RVT U3454 ( .A(\u_div/SumTmp[20][0] ), .Y(net31203) );
  INVX0_RVT U3455 ( .A(\u_div/SumTmp[10][9] ), .Y(net31204) );
  INVX0_RVT U3456 ( .A(\u_div/SumTmp[11][8] ), .Y(net31205) );
  INVX0_RVT U3457 ( .A(\u_div/SumTmp[12][7] ), .Y(net31206) );
  INVX0_RVT U3458 ( .A(\u_div/SumTmp[13][6] ), .Y(net31207) );
  INVX0_RVT U3459 ( .A(\u_div/SumTmp[14][5] ), .Y(net31208) );
  INVX0_RVT U3460 ( .A(\u_div/SumTmp[15][4] ), .Y(net31209) );
  INVX0_RVT U3461 ( .A(\u_div/SumTmp[17][2] ), .Y(net31211) );
  INVX0_RVT U3462 ( .A(\u_div/SumTmp[18][1] ), .Y(net31212) );
  INVX0_RVT U3463 ( .A(\u_div/SumTmp[19][0] ), .Y(net31213) );
  AND2X1_RVT U3464 ( .A1(n1203), .A2(net37169), .Y(quotient[46]) );
  AND4X1_RVT U3465 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .Y(n1203)
         );
  NOR3X0_RVT U3466 ( .A1(net32210), .A2(net32300), .A3(net32324), .Y(n1207) );
  NOR2X0_RVT U3467 ( .A1(net32264), .A2(net32234), .Y(n1206) );
  NOR2X0_RVT U3468 ( .A1(b[1]), .A2(b[2]), .Y(n1205) );
  NOR2X0_RVT U3469 ( .A1(net32352), .A2(n1014), .Y(n1204) );
  NOR2X0_RVT U3470 ( .A1(n1208), .A2(n1209), .Y(quotient[45]) );
  NAND4X0_RVT U3471 ( .A1(n1210), .A2(n1211), .A3(n1212), .A4(n1213), .Y(n1209) );
  NOR3X0_RVT U3472 ( .A1(net32234), .A2(net32210), .A3(net32178), .Y(n1213) );
  NOR3X0_RVT U3473 ( .A1(net32300), .A2(net32264), .A3(net32324), .Y(n1212) );
  NOR3X0_RVT U3474 ( .A1(b[2]), .A2(net31814), .A3(net32352), .Y(n1211) );
  NOR3X0_RVT U3475 ( .A1(net31872), .A2(net31896), .A3(net31844), .Y(n1210) );
  NAND4X0_RVT U3476 ( .A1(n1214), .A2(n1215), .A3(n1216), .A4(n1217), .Y(n1208) );
  NOR3X0_RVT U3477 ( .A1(net31950), .A2(net31972), .A3(net31922), .Y(n1217) );
  NOR3X0_RVT U3478 ( .A1(net32024), .A2(b[14]), .A3(net31998), .Y(n1216) );
  NOR3X0_RVT U3479 ( .A1(net32104), .A2(net32128), .A3(net32076), .Y(n1215) );
  NOR2X0_RVT U3480 ( .A1(net32154), .A2(n1114), .Y(n1214) );
  NAND4X0_RVT U3481 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .Y(
        net31244) );
  NOR3X0_RVT U3482 ( .A1(net32234), .A2(net32210), .A3(net32178), .Y(n1221) );
  NOR3X0_RVT U3483 ( .A1(net32300), .A2(net32264), .A3(net32324), .Y(n1220) );
  NOR3X0_RVT U3484 ( .A1(net31844), .A2(net31814), .A3(net31872), .Y(n1219) );
  NOR2X0_RVT U3485 ( .A1(net31896), .A2(net31922), .Y(n1218) );
  NAND4X0_RVT U3486 ( .A1(net32046), .A2(net32016), .A3(net31986), .A4(n1222), 
        .Y(net31242) );
  NAND4X0_RVT U3487 ( .A1(\u_div/CryTmp[42][5] ), .A2(n1224), .A3(n1225), .A4(
        n1226), .Y(n1223) );
  NOR2X0_RVT U3488 ( .A1(net32178), .A2(net32210), .Y(n1226) );
  NOR2X0_RVT U3489 ( .A1(net32234), .A2(net32264), .Y(n1225) );
  NOR2X0_RVT U3490 ( .A1(net32300), .A2(net32154), .Y(n1224) );
  NAND4X0_RVT U3491 ( .A1(\u_div/CryTmp[41][6] ), .A2(net32156), .A3(n1227), 
        .A4(n1228), .Y(net31261) );
  NOR2X0_RVT U3492 ( .A1(net32178), .A2(net32210), .Y(n1228) );
  NOR2X0_RVT U3493 ( .A1(net32234), .A2(net32264), .Y(n1227) );
  NAND2X0_RVT U3494 ( .A1(\u_div/CryTmp[40][7] ), .A2(net32156), .Y(n1230) );
  NAND2X0_RVT U3495 ( .A1(net32226), .A2(net32186), .Y(n1229) );
  AND2X1_RVT U3496 ( .A1(n1231), .A2(n1232), .Y(net31273) );
  NOR3X0_RVT U3497 ( .A1(net31950), .A2(net32178), .A3(net31922), .Y(n1232) );
  NOR3X0_RVT U3498 ( .A1(net32024), .A2(net31972), .A3(net31998), .Y(n1231) );
  NOR3X0_RVT U3499 ( .A1(net32104), .A2(b[14]), .A3(net32076), .Y(net31271) );
  NOR2X0_RVT U3500 ( .A1(net32128), .A2(net32154), .Y(net31270) );
  NAND4X0_RVT U3501 ( .A1(n1233), .A2(n1234), .A3(n1235), .A4(n1236), .Y(
        net31255) );
  NOR4X0_RVT U3502 ( .A1(net31814), .A2(net31844), .A3(net31872), .A4(net31896), .Y(n1236) );
  NOR3X0_RVT U3503 ( .A1(net31972), .A2(net31922), .A3(net31950), .Y(n1235) );
  NOR3X0_RVT U3504 ( .A1(b[14]), .A2(net31998), .A3(net32024), .Y(n1234) );
  NOR3X0_RVT U3505 ( .A1(net32128), .A2(net32076), .A3(net32104), .Y(n1233) );
  OR2X1_RVT U3506 ( .A1(net32076), .A2(net31292), .Y(net31287) );
  OR4X1_RVT U3507 ( .A1(net32024), .A2(b[14]), .A3(net31998), .A4(net31295), 
        .Y(net31292) );
  OR3X1_RVT U3508 ( .A1(n1237), .A2(n1238), .A3(n1239), .Y(net31295) );
  OR3X1_RVT U3509 ( .A1(net31922), .A2(net31950), .A3(net31972), .Y(n1239) );
  OR2X1_RVT U3510 ( .A1(net31872), .A2(net31896), .Y(n1238) );
  OR2X1_RVT U3511 ( .A1(net31814), .A2(net31844), .Y(n1237) );
  OR4X1_RVT U3512 ( .A1(net31844), .A2(net31814), .A3(net31896), .A4(net31872), 
        .Y(net31276) );
endmodule


module fpu ( clk, rst, a, b, sel, err, overflow, y );
  input [31:0] a;
  input [31:0] b;
  input [1:0] sel;
  output [31:0] y;
  input clk, rst;
  output err, overflow;
  wire   tmp_s0, tmp_a_s1, tmp_b_s1, \sel_2[1] , N94, N95, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N255, N256, N257, N258, N350, N351, N352, N353, N354, N355, N356,
         N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367,
         N368, N369, N370, N371, N372, N373, N374, N408, N409, N410, N411,
         N412, N413, N414, N415, N416, N417, N418, N419, N420, N421, N422,
         N423, N424, N425, N426, N427, N428, N429, N430, N431, N432, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445,
         N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
         N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467,
         N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478,
         N479, N480, N481, N482, N483, N928, N929, N930, N931, N932, N933,
         N934, N935, N936, N937, N938, N939, N940, N941, N942, N943, N944,
         N945, N946, N947, N948, N949, N950, N951, N952, N953, N954, N955,
         N956, N957, N958, N959, N960, N961, N962, N963, N964, N965, N966,
         N967, N968, N969, N970, N971, N972, N973, N974, N975, N976, N977,
         N978, N979, N980, N981, N982, N983, N984, N993, N994, N995, N996,
         N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006,
         N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016,
         N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026,
         N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036,
         N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046,
         N1047, N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056,
         N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066,
         N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076,
         N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086,
         N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096,
         N1097, N1098, N1099, N1116, N1117, N1118, N1119, N1120, N1121, N1122,
         N1123, N1124, N1129, N1131, N1132, N1133, N1134, N1135, N1136, N1137,
         N1138, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148,
         N1188, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1198, N1199,
         N1200, N1201, N1202, N1203, N1204, N1205, N1206, N1249, N1250, N1251,
         N1252, N1253, N1254, N1255, N1256, N1258, N1259, N1260, N1261, N1262,
         N1263, N1264, N1265, N1266, N1314, N1315, N1316, N1317, N1318, N1320,
         N1321, N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1382, N1383,
         N1384, N1385, N1386, N1387, N1388, N1389, N1391, N1392, N1393, N1394,
         N1395, N1396, N1397, N1398, N1399, N1449, N1450, N1451, N1452, N1453,
         N1454, N1455, N1457, N1458, N1459, N1460, N1461, N1462, N1463, N1464,
         N1465, N1516, N1517, N1518, N1519, N1520, N1521, N1522, N1523, N1525,
         N1526, N1527, N1528, N1529, N1530, N1531, N1532, N1533, N1588, N1589,
         N1590, N1591, N1592, N1593, N1595, N1596, N1597, N1598, N1599, N1600,
         N1601, N1602, N1603, N1661, N1662, N1663, N1664, N1665, N1666, N1667,
         N1668, N1670, N1671, N1672, N1673, N1674, N1675, N1676, N1677, N1678,
         N1736, N1737, N1738, N1739, N1740, N1741, N1742, N1744, N1745, N1746,
         N1747, N1748, N1749, N1750, N1751, N1752, N1811, N1812, N1813, N1814,
         N1815, N1816, N1817, N1818, N1820, N1821, N1822, N1823, N1824, N1825,
         N1826, N1827, N1828, N1886, N1887, N1888, N1889, N1890, N1891, N1892,
         N1893, N1894, N1895, N1958, N1959, N1960, N1961, N1962, N1963, N1964,
         N1965, N1967, N1968, N1969, N1970, N1971, N1972, N1973, N1974, N1975,
         N2036, N2037, N2038, N2039, N2040, N2041, N2042, N2043, N2044, N2047,
         N2048, N2049, N2050, N2051, N2052, N2053, N2054, N2055, N2056, N2057,
         N2058, N2059, N2060, N2061, N2062, N2063, N2064, N2065, N2066, N2067,
         N2068, N2069, N2070, N2071, N2072, N2073, N2074, N2078, N2079, N2080,
         N2081, N2084, N2085, N2086, N2087, N2088, N2089, N2090, N2091, N2092,
         N2093, N2094, N2095, N2096, N2097, N2098, N2099, N2100, N2101, N2102,
         N2103, N2104, N2105, N2106, N2107, N2108, N2109, N2110, N2111, N2112,
         N2118, N2119, N2131, N2132, N2206, N2207, N2208, N2209, N2210, N2211,
         N2212, N2213, N2214, N2215, N2216, N2217, N2218, N2219, N2220, N2221,
         N2222, N2223, N2224, N2225, N2226, N2227, N2228, N2230, N2233, N2235,
         N2236, N2237, N2238, N2239, N2240, N2241, N2242, N2243, N2244, N2245,
         N2246, N2247, N2248, N2249, N2250, N2251, N2252, N2253, N2254, N2255,
         N2256, N2257, N2258, N2259, N2260, N2261, N2262, N2263, N2264, N2295,
         N2296, N2297, N2298, N2299, N2300, N2301, N2302, N2303, N2304, N2305,
         N2306, N2307, N2308, N2309, N2310, N2311, N2312, N2313, N2314, N2315,
         N2316, N2450, N2463, N2464, N2465, N2466, N2467, N2468, N2469, N2470,
         N2471, N2472, N2473, N2474, N2475, N2476, N2477, N2478, N2479, N2480,
         N2481, N2482, N2483, N2484, N2515, N2516, N2517, N2518, N2519, N2520,
         N2521, N2522, N2523, N2524, N2525, N2526, N2527, N2528, N2529, N2530,
         N2531, N2532, N2533, N2534, N2535, N2536, N2768, N2769, N2770, N2771,
         N2772, N2773, N2774, N2775, N2776, N2777, N2778, N2779, N2780, N2781,
         N2782, N2783, N2784, N2785, N2786, N2787, N2788, N2789, N2790, N2791,
         N2792, N2793, N2794, N2795, N2796, N2797, N2798, N2799, N2800, N2801,
         n153, n154, n156, n157, n158, n159, n161, n163, n164, n166, n167,
         n168, n169, n172, n173, n175, n176, n177, n178, n180, n181, n184,
         n185, n186, n189, n190, n193, n194, n197, n198, n201, n202, n205,
         n206, n209, n210, n213, n214, n218, n220, n221, n223, n224, n225,
         n226, n228, n229, n230, n231, n232, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n330,
         n333, n334, n339, n340, n342, n343, n344, n345, n346, n347, n349,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n366, n367, n368, n369, n370, n371, n372, n373, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n386, n389, n390, n391, n392,
         n398, n399, n400, n401, n402, n408, n418, n419, n420, n421, n426,
         n428, n432, n452, n454, n455, n456, n457, n458, n459, n461, n462,
         n463, n464, n466, n467, n470, n471, n472, n473, n475, n479, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n553, n555, n556, n557,
         n558, n559, n560, n561, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n573, n574, n576, n577, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n625, n626, n627, n628, n629, n630,
         n634, n635, n636, n643, n644, n647, n648, n849, n850, n851, n855,
         n856, n857, n858, n867, n869, n870, n871, n879, n880, n883, n884,
         n885, n886, n887, n892, n893, n896, n897, n898, n899, n900, n905,
         n906, n909, n910, n911, n912, n913, n918, n919, n922, n923, n924,
         n925, n926, n931, n932, n935, n936, n937, n938, n939, n944, n945,
         n948, n949, n950, n951, n952, n957, n958, n961, n962, n963, n964,
         n965, n967, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n984, n987, n988, n989, n990, n991, n994,
         n1000, n1002, n1005, n1006, n1007, n1015, n1031, n1136, n1137, n1138,
         n1139, n1140, n1141, n1143, n1144, n1147, n1148, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1174,
         n1175, n1176, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1190, n1192, n1194, n1196, n1198, n1200, n1202,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1254, n1255,
         n1256, n1257, n1258, n1260, n1261, n1262, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, \add_489/carry[8] , \add_489/carry[7] , \add_489/carry[6] ,
         \add_489/carry[5] , \add_489/carry[4] , \add_489/carry[3] ,
         \add_480/carry[2] , \add_480/carry[3] , \add_480/carry[4] ,
         \add_480/carry[5] , \add_480/carry[6] , \add_480/carry[7] ,
         \add_480/carry[8] , \add_480/carry[9] , \sub_467/carry[2] ,
         \sub_467/carry[3] , \sub_467/carry[4] , \sub_467/carry[5] ,
         \sub_467/carry[6] , \sub_467/carry[7] , \sub_467/carry[8] ,
         \sub_467/carry[9] , \sub_458/carry[9] , \sub_458/carry[8] ,
         \sub_458/carry[7] , \sub_458/carry[6] , \sub_458/carry[5] ,
         \sub_458/carry[4] , \sub_458/carry[3] , \sub_424/carry[9] ,
         \sub_424/carry[8] , \sub_424/carry[7] , \sub_424/carry[6] ,
         \sub_424/carry[5] , \sub_424/carry[4] , \sub_424/carry[3] ,
         \sub_413/carry[2] , \sub_413/carry[3] , \sub_413/carry[4] ,
         \sub_413/carry[5] , \sub_413/carry[6] , \sub_413/carry[7] ,
         \sub_413/carry[8] , \sub_413/carry[9] , \sub_408/carry[9] ,
         \sub_408/carry[8] , \sub_408/carry[7] , \sub_408/carry[6] ,
         \sub_408/carry[5] , \sub_408/carry[4] , \sub_400/carry[2] ,
         \sub_400/carry[3] , \sub_400/carry[4] , \sub_400/carry[5] ,
         \sub_400/carry[6] , \sub_400/carry[7] , \sub_400/carry[8] ,
         \sub_400/carry[9] , \sub_395/carry[9] , \sub_395/carry[8] ,
         \sub_395/carry[7] , \sub_395/carry[6] , \sub_395/carry[5] ,
         \sub_395/carry[4] , \sub_395/carry[3] , \sub_381/carry[2] ,
         \sub_381/carry[3] , \sub_381/carry[4] , \sub_381/carry[5] ,
         \sub_381/carry[6] , \sub_381/carry[7] , \sub_381/carry[8] ,
         \sub_381/carry[9] , \sub_376/carry[9] , \sub_376/carry[8] ,
         \sub_376/carry[7] , \sub_376/carry[6] , \sub_376/carry[5] ,
         \sub_368/carry[2] , \sub_368/carry[3] , \sub_368/carry[4] ,
         \sub_368/carry[5] , \sub_368/carry[6] , \sub_368/carry[7] ,
         \sub_368/carry[8] , \sub_368/carry[9] , \sub_363/carry[9] ,
         \sub_363/carry[8] , \sub_363/carry[7] , \sub_363/carry[6] ,
         \sub_363/carry[5] , \sub_363/carry[4] , \sub_363/carry[3] ,
         \sub_352/carry[2] , \sub_352/carry[3] , \sub_352/carry[4] ,
         \sub_352/carry[5] , \sub_352/carry[6] , \sub_352/carry[7] ,
         \sub_352/carry[8] , \sub_352/carry[9] , \sub_347/carry[9] ,
         \sub_347/carry[8] , \sub_347/carry[7] , \sub_347/carry[6] ,
         \sub_347/carry[5] , \sub_347/carry[4] , \sub_339/carry[2] ,
         \sub_339/carry[3] , \sub_339/carry[4] , \sub_339/carry[5] ,
         \sub_339/carry[6] , \sub_339/carry[7] , \sub_339/carry[8] ,
         \sub_339/carry[9] , \sub_334/carry[9] , \sub_334/carry[8] ,
         \sub_334/carry[7] , \sub_334/carry[6] , \sub_334/carry[5] ,
         \sub_334/carry[4] , \sub_334/carry[3] , \sub_317/carry[2] ,
         \sub_317/carry[3] , \sub_317/carry[4] , \sub_317/carry[5] ,
         \sub_317/carry[6] , \sub_317/carry[7] , \sub_317/carry[8] ,
         \sub_317/carry[9] , \sub_312/carry[9] , \sub_312/carry[8] ,
         \sub_312/carry[7] , \sub_312/carry[6] , \sub_304/carry[2] ,
         \sub_304/carry[3] , \sub_304/carry[4] , \sub_304/carry[5] ,
         \sub_304/carry[6] , \sub_304/carry[7] , \sub_304/carry[8] ,
         \sub_304/carry[9] , \sub_299/carry[9] , \sub_299/carry[8] ,
         \sub_299/carry[7] , \sub_299/carry[6] , \sub_299/carry[5] ,
         \sub_299/carry[4] , \sub_299/carry[3] , \sub_288/carry[2] ,
         \sub_288/carry[3] , \sub_288/carry[4] , \sub_288/carry[5] ,
         \sub_288/carry[6] , \sub_288/carry[7] , \sub_288/carry[8] ,
         \sub_288/carry[9] , \sub_283/carry[9] , \sub_283/carry[8] ,
         \sub_283/carry[7] , \sub_283/carry[6] , \sub_283/carry[5] ,
         \sub_283/carry[4] , \sub_275/carry[2] , \sub_275/carry[3] ,
         \sub_275/carry[4] , \sub_275/carry[5] , \sub_275/carry[6] ,
         \sub_275/carry[7] , \sub_275/carry[8] , \sub_275/carry[9] ,
         \sub_270/carry[9] , \sub_270/carry[8] , \sub_270/carry[7] ,
         \sub_270/carry[6] , \sub_270/carry[5] , \sub_270/carry[4] ,
         \sub_270/carry[3] , \sub_259/carry[2] , \sub_259/carry[3] ,
         \sub_259/carry[4] , \sub_259/carry[5] , \sub_259/carry[6] ,
         \sub_259/carry[7] , \sub_259/carry[8] , \sub_259/carry[9] , net27434,
         net27435, net27438, net27580, net27586, net32870, net32868, net32866,
         net32864, net32882, net32880, net32878, net32876, net32926, net32924,
         net32932, net32930, net32938, net32948, net32946, net32952, net32950,
         net32958, net32956, net32962, net36423, net47575, net47581, net47614,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487;
  wire   [7:0] a_e;
  wire   [23:0] a_m;
  wire   [7:0] b_e;
  wire   [23:0] b_m;
  wire   [1:0] sel_0;
  wire   [1:0] sel_1;
  wire   [47:0] tmp_m0;
  wire   [7:0] tmp_a_e1;
  wire   [22:0] tmp_a_m1;
  wire   [7:0] tmp_b_e1;
  wire   [22:0] tmp_b_m1;
  wire   [9:0] tmp_e1;
  wire   [47:0] tmp_m1;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23;

  DFFARX1_RVT \tmp_m1_reg[23]  ( .D(N2088), .CLK(clk), .RSTB(n1975), .Q(
        tmp_m1[23]) );
  DFFARX1_RVT \tmp_m1_reg[0]  ( .D(N2065), .CLK(clk), .RSTB(n1975), .Q(
        tmp_m1[0]), .QN(n1617) );
  AOI21X1_RVT U138 ( .A1(n164), .A2(n2445), .A3(n166), .Y(n163) );
  NAND2X0_RVT U141 ( .A1(n2443), .A2(n172), .Y(n168) );
  NAND3X0_RVT U145 ( .A1(n176), .A2(n177), .A3(n178), .Y(N2799) );
  NAND2X0_RVT U147 ( .A1(N2242), .A2(n184), .Y(n177) );
  NAND3X0_RVT U148 ( .A1(n176), .A2(n185), .A3(n186), .Y(N2798) );
  NAND2X0_RVT U150 ( .A1(N2241), .A2(n184), .Y(n185) );
  NAND3X0_RVT U151 ( .A1(n176), .A2(n189), .A3(n190), .Y(N2797) );
  NAND2X0_RVT U153 ( .A1(N2240), .A2(n184), .Y(n189) );
  NAND3X0_RVT U154 ( .A1(n176), .A2(n193), .A3(n194), .Y(N2796) );
  NAND2X0_RVT U156 ( .A1(N2239), .A2(n184), .Y(n193) );
  NAND3X0_RVT U157 ( .A1(n176), .A2(n197), .A3(n198), .Y(N2795) );
  NAND2X0_RVT U159 ( .A1(N2238), .A2(n184), .Y(n197) );
  NAND3X0_RVT U160 ( .A1(n176), .A2(n201), .A3(n202), .Y(N2794) );
  NAND2X0_RVT U164 ( .A1(N2237), .A2(n184), .Y(n201) );
  NAND3X0_RVT U165 ( .A1(n176), .A2(n205), .A3(n206), .Y(N2793) );
  NAND2X0_RVT U169 ( .A1(N2236), .A2(n184), .Y(n205) );
  NAND3X0_RVT U170 ( .A1(n176), .A2(n209), .A3(n210), .Y(N2792) );
  NOR4X0_RVT U173 ( .A1(n213), .A2(n214), .A3(n1832), .A4(n1841), .Y(n181) );
  NAND2X0_RVT U175 ( .A1(N2235), .A2(n184), .Y(n209) );
  NAND3X0_RVT U178 ( .A1(n224), .A2(n225), .A3(n226), .Y(n220) );
  NAND2X0_RVT U179 ( .A1(n2450), .A2(n228), .Y(n218) );
  AND3X1_RVT U186 ( .A1(n238), .A2(n239), .A3(\sel_2[1] ), .Y(n223) );
  NAND3X0_RVT U187 ( .A1(n240), .A2(n172), .A3(n226), .Y(n238) );
  NAND2X0_RVT U188 ( .A1(n241), .A2(n242), .Y(n240) );
  OAI221X1_RVT U190 ( .A1(n172), .A2(n224), .A3(n242), .A4(n225), .A5(n226), 
        .Y(n237) );
  NAND2X0_RVT U304 ( .A1(n333), .A2(n334), .Y(n213) );
  NAND4X0_RVT U305 ( .A1(n2445), .A2(n2448), .A3(n239), .A4(n1617), .Y(n334)
         );
  NAND4X0_RVT U306 ( .A1(n2445), .A2(n164), .A3(n2474), .A4(n1617), .Y(n333)
         );
  NAND3X0_RVT U315 ( .A1(n345), .A2(n172), .A3(n2448), .Y(n344) );
  NAND2X0_RVT U318 ( .A1(n226), .A2(n2449), .Y(n224) );
  NAND2X0_RVT U319 ( .A1(n226), .A2(n2465), .Y(n225) );
  AND3X1_RVT U321 ( .A1(n2445), .A2(n349), .A3(tmp_m1[0]), .Y(n328) );
  NAND2X0_RVT U324 ( .A1(n226), .A2(\sel_2[1] ), .Y(n156) );
  AND3X1_RVT U325 ( .A1(n2445), .A2(n2475), .A3(tmp_m1[23]), .Y(n330) );
  NAND2X0_RVT U327 ( .A1(\sel_2[1] ), .A2(n2476), .Y(n239) );
  NAND4X0_RVT U329 ( .A1(n347), .A2(n2450), .A3(n2485), .A4(n2486), .Y(n157)
         );
  NAND3X0_RVT U333 ( .A1(n2443), .A2(n2474), .A3(n2441), .Y(n180) );
  NAND2X0_RVT U338 ( .A1(n228), .A2(n353), .Y(n166) );
  NAND3X0_RVT U339 ( .A1(n347), .A2(n164), .A3(n346), .Y(n353) );
  AND3X1_RVT U340 ( .A1(n2450), .A2(n2485), .A3(N2119), .Y(n346) );
  NAND2X0_RVT U342 ( .A1(n2444), .A2(n164), .Y(n228) );
  NAND3X0_RVT U344 ( .A1(n347), .A2(n2450), .A3(N2118), .Y(n343) );
  NAND4X0_RVT U346 ( .A1(n2469), .A2(n2468), .A3(n354), .A4(n355), .Y(n172) );
  NOR4X0_RVT U347 ( .A1(n356), .A2(tmp_b_e1[0]), .A3(tmp_b_e1[1]), .A4(
        tmp_b_e1[2]), .Y(n355) );
  AND3X1_RVT U348 ( .A1(n2466), .A2(n2464), .A3(n2467), .Y(n354) );
  NAND4X0_RVT U354 ( .A1(n2454), .A2(n2453), .A3(n357), .A4(n358), .Y(n242) );
  NOR4X0_RVT U355 ( .A1(n359), .A2(tmp_a_e1[0]), .A3(tmp_a_e1[1]), .A4(
        tmp_a_e1[2]), .Y(n358) );
  AND3X1_RVT U356 ( .A1(n2451), .A2(n2446), .A3(n2452), .Y(n357) );
  NAND2X0_RVT U362 ( .A1(n2450), .A2(n164), .Y(n167) );
  NAND3X0_RVT U363 ( .A1(N2131), .A2(n360), .A3(N2132), .Y(n164) );
  XNOR3X1_RVT U364 ( .A1(tmp_b_s1), .A2(tmp_a_s1), .A3(n2476), .Y(n360) );
  NAND2X0_RVT U367 ( .A1(n175), .A2(n169), .Y(n241) );
  AOI22X1_RVT U369 ( .A1(n2449), .A2(n359), .A3(n2465), .A4(n356), .Y(n226) );
  NAND4X0_RVT U371 ( .A1(n2460), .A2(n2459), .A3(n366), .A4(n367), .Y(n363) );
  NOR4X0_RVT U372 ( .A1(tmp_b_m1[15]), .A2(tmp_b_m1[16]), .A3(tmp_b_m1[14]), 
        .A4(n368), .Y(n367) );
  NOR3X0_RVT U374 ( .A1(tmp_b_m1[12]), .A2(tmp_b_m1[13]), .A3(tmp_b_m1[11]), 
        .Y(n366) );
  OR4X1_RVT U377 ( .A1(tmp_b_m1[20]), .A2(tmp_b_m1[21]), .A3(tmp_b_m1[1]), 
        .A4(n369), .Y(n362) );
  OR4X1_RVT U379 ( .A1(tmp_b_m1[5]), .A2(tmp_b_m1[6]), .A3(tmp_b_m1[4]), .A4(
        n370), .Y(n361) );
  NAND4X0_RVT U383 ( .A1(n2463), .A2(n2462), .A3(n376), .A4(n377), .Y(n373) );
  NOR4X0_RVT U384 ( .A1(tmp_a_m1[15]), .A2(tmp_a_m1[16]), .A3(tmp_a_m1[14]), 
        .A4(n378), .Y(n377) );
  NOR3X0_RVT U386 ( .A1(tmp_a_m1[12]), .A2(tmp_a_m1[13]), .A3(tmp_a_m1[11]), 
        .Y(n376) );
  OR4X1_RVT U389 ( .A1(tmp_a_m1[20]), .A2(tmp_a_m1[21]), .A3(tmp_a_m1[1]), 
        .A4(n379), .Y(n372) );
  OR4X1_RVT U391 ( .A1(tmp_a_m1[5]), .A2(tmp_a_m1[6]), .A3(tmp_a_m1[4]), .A4(
        n380), .Y(n371) );
  NAND4X0_RVT U395 ( .A1(tmp_b_e1[7]), .A2(tmp_b_e1[6]), .A3(tmp_b_e1[5]), 
        .A4(tmp_b_e1[4]), .Y(n382) );
  NAND4X0_RVT U396 ( .A1(tmp_b_e1[3]), .A2(tmp_b_e1[2]), .A3(tmp_b_e1[1]), 
        .A4(tmp_b_e1[0]), .Y(n381) );
  NAND4X0_RVT U398 ( .A1(tmp_a_e1[7]), .A2(tmp_a_e1[6]), .A3(tmp_a_e1[5]), 
        .A4(tmp_a_e1[4]), .Y(n384) );
  NAND4X0_RVT U399 ( .A1(tmp_a_e1[3]), .A2(tmp_a_e1[2]), .A3(tmp_a_e1[1]), 
        .A4(tmp_a_e1[0]), .Y(n383) );
  NAND4X0_RVT U401 ( .A1(n389), .A2(n390), .A3(n391), .A4(n392), .Y(n386) );
  NAND2X0_RVT U418 ( .A1(n454), .A2(n455), .Y(n452) );
  NAND4X0_RVT U424 ( .A1(n470), .A2(n471), .A3(n472), .A4(n473), .Y(n466) );
  NAND4X0_RVT U440 ( .A1(n490), .A2(n491), .A3(n492), .A4(n493), .Y(n488) );
  NAND4X0_RVT U455 ( .A1(n504), .A2(n505), .A3(n506), .A4(n507), .Y(n503) );
  AOI222X1_RVT U469 ( .A1(n1901), .A2(tmp_m0[39]), .A3(n2320), .A4(n518), .A5(
        n1863), .A6(tmp_m0[40]), .Y(n513) );
  NAND4X0_RVT U470 ( .A1(n519), .A2(n520), .A3(n521), .A4(n522), .Y(n518) );
  AOI222X1_RVT U482 ( .A1(n1901), .A2(tmp_m0[38]), .A3(n2320), .A4(n529), .A5(
        n1863), .A6(tmp_m0[39]), .Y(n527) );
  NAND4X0_RVT U483 ( .A1(n530), .A2(n531), .A3(n532), .A4(n533), .Y(n529) );
  NAND4X0_RVT U519 ( .A1(n558), .A2(n559), .A3(n560), .A4(n561), .Y(n556) );
  NAND4X0_RVT U543 ( .A1(n585), .A2(n586), .A3(n587), .A4(n588), .Y(n583) );
  NAND4X0_RVT U553 ( .A1(n593), .A2(n594), .A3(n595), .A4(n596), .Y(n591) );
  NAND4X0_RVT U562 ( .A1(n600), .A2(n601), .A3(n602), .A4(n603), .Y(n598) );
  NAND4X0_RVT U570 ( .A1(n606), .A2(n607), .A3(n608), .A4(n609), .Y(n604) );
  NAND4X0_RVT U578 ( .A1(n612), .A2(n613), .A3(n614), .A4(n615), .Y(n610) );
  NAND4X0_RVT U592 ( .A1(n628), .A2(n626), .A3(n627), .A4(n625), .Y(n623) );
  AND3X1_RVT U624 ( .A1(n647), .A2(n648), .A3(n1894), .Y(n643) );
  NAND2X0_RVT U944 ( .A1(n972), .A2(n973), .Y(n971) );
  NOR4X0_RVT U945 ( .A1(n974), .A2(n975), .A3(n976), .A4(n977), .Y(n973) );
  NAND2X0_RVT U961 ( .A1(n2473), .A2(n1561), .Y(n849) );
  NOR4X0_RVT U969 ( .A1(n988), .A2(n989), .A3(n990), .A4(n991), .Y(n987) );
  NAND2X0_RVT U1247 ( .A1(n1140), .A2(n1143), .Y(n1144) );
  NAND2X0_RVT U1255 ( .A1(n1153), .A2(n1154), .Y(n1152) );
  AND3X1_RVT U1257 ( .A1(n1609), .A2(n2325), .A3(n1158), .Y(n1157) );
  NAND4X0_RVT U1259 ( .A1(n2437), .A2(n1160), .A3(n1161), .A4(n1137), .Y(n1156) );
  NAND2X0_RVT U1260 ( .A1(sel_0[0]), .A2(n2440), .Y(n1137) );
  NAND2X0_RVT U1262 ( .A1(sel_0[0]), .A2(n2323), .Y(n1161) );
  NAND2X0_RVT U1264 ( .A1(n2326), .A2(n2325), .Y(n1160) );
  NAND2X0_RVT U1300 ( .A1(n1150), .A2(n1148), .Y(n1162) );
  NAND2X0_RVT U1302 ( .A1(N95), .A2(n2439), .Y(n1150) );
  NAND2X0_RVT U1307 ( .A1(n1138), .A2(n1140), .Y(n1158) );
  NAND2X0_RVT U1309 ( .A1(N94), .A2(n1147), .Y(n1138) );
  AOI21X1_RVT U1310 ( .A1(n1136), .A2(n1176), .A3(sel_0[0]), .Y(n1175) );
  NAND2X0_RVT U1311 ( .A1(n2326), .A2(N94), .Y(n1136) );
  NAND2X0_RVT U1312 ( .A1(n1141), .A2(n1139), .Y(n1155) );
  NAND2X0_RVT U1313 ( .A1(n1781), .A2(N94), .Y(n1139) );
  NAND2X0_RVT U1314 ( .A1(n1781), .A2(n2324), .Y(n1141) );
  OR3X2_RVT U180 ( .A1(n229), .A2(n230), .A3(n231), .Y(N2791) );
  OR3X2_RVT U191 ( .A1(n244), .A2(n245), .A3(n246), .Y(N2790) );
  OR3X2_RVT U196 ( .A1(n248), .A2(n249), .A3(n250), .Y(N2789) );
  OR3X2_RVT U201 ( .A1(n252), .A2(n253), .A3(n254), .Y(N2788) );
  OR3X2_RVT U206 ( .A1(n256), .A2(n257), .A3(n258), .Y(N2787) );
  OR3X2_RVT U211 ( .A1(n260), .A2(n261), .A3(n262), .Y(N2786) );
  OR3X2_RVT U216 ( .A1(n264), .A2(n265), .A3(n266), .Y(N2785) );
  OR3X2_RVT U221 ( .A1(n268), .A2(n269), .A3(n270), .Y(N2784) );
  OR3X2_RVT U226 ( .A1(n272), .A2(n273), .A3(n274), .Y(N2783) );
  OR3X2_RVT U231 ( .A1(n276), .A2(n277), .A3(n278), .Y(N2782) );
  OR3X2_RVT U236 ( .A1(n280), .A2(n281), .A3(n282), .Y(N2781) );
  OR3X2_RVT U241 ( .A1(n284), .A2(n285), .A3(n286), .Y(N2780) );
  OR3X2_RVT U246 ( .A1(n288), .A2(n289), .A3(n290), .Y(N2779) );
  OR3X2_RVT U251 ( .A1(n292), .A2(n293), .A3(n294), .Y(N2778) );
  OR3X2_RVT U256 ( .A1(n296), .A2(n297), .A3(n298), .Y(N2777) );
  OR3X2_RVT U261 ( .A1(n300), .A2(n301), .A3(n302), .Y(N2776) );
  OR3X2_RVT U266 ( .A1(n304), .A2(n305), .A3(n306), .Y(N2775) );
  OR3X2_RVT U271 ( .A1(n308), .A2(n309), .A3(n310), .Y(N2774) );
  OR3X2_RVT U276 ( .A1(n312), .A2(n313), .A3(n314), .Y(N2773) );
  OR3X2_RVT U281 ( .A1(n316), .A2(n317), .A3(n318), .Y(N2772) );
  OR3X2_RVT U286 ( .A1(n320), .A2(n321), .A3(n322), .Y(N2771) );
  OR3X2_RVT U291 ( .A1(n324), .A2(n325), .A3(n326), .Y(N2770) );
  OR3X2_RVT U370 ( .A1(n361), .A2(n362), .A3(n363), .Y(n356) );
  OR3X2_RVT U373 ( .A1(tmp_b_m1[18]), .A2(tmp_b_m1[19]), .A3(tmp_b_m1[17]), 
        .Y(n368) );
  OR3X2_RVT U378 ( .A1(tmp_b_m1[2]), .A2(tmp_b_m1[3]), .A3(tmp_b_m1[22]), .Y(
        n369) );
  OR3X2_RVT U380 ( .A1(tmp_b_m1[8]), .A2(tmp_b_m1[9]), .A3(tmp_b_m1[7]), .Y(
        n370) );
  OR3X2_RVT U382 ( .A1(n371), .A2(n372), .A3(n373), .Y(n359) );
  OR3X2_RVT U385 ( .A1(tmp_a_m1[18]), .A2(tmp_a_m1[19]), .A3(tmp_a_m1[17]), 
        .Y(n378) );
  OR3X2_RVT U390 ( .A1(tmp_a_m1[2]), .A2(tmp_a_m1[3]), .A3(tmp_a_m1[22]), .Y(
        n379) );
  OR3X2_RVT U392 ( .A1(tmp_a_m1[8]), .A2(tmp_a_m1[9]), .A3(tmp_a_m1[7]), .Y(
        n380) );
  OR3X2_RVT U1306 ( .A1(n1155), .A2(n1175), .A3(n1158), .Y(n1174) );
  fpu_DW01_inc_0 add_706 ( .A(tmp_m1[45:24]), .SUM({N2536, N2535, N2534, N2533, 
        N2532, N2531, N2530, N2529, N2528, N2527, N2526, N2525, N2524, N2523, 
        N2522, N2521, N2520, N2519, N2518, N2517, N2516, N2515}) );
  fpu_DW01_inc_1 add_699_2 ( .A(tmp_m1[46:25]), .SUM({N2484, N2483, N2482, 
        N2481, N2480, N2479, N2478, N2477, N2476, N2475, N2474, N2473, N2472, 
        N2471, N2470, N2469, N2468, N2467, N2466, N2465, N2464, N2463}) );
  fpu_DW01_inc_2 add_442 ( .A({n1927, n1923, n1921, n1919, n1917, n1913, n1902, 
        n1906, n1909, n1911}), .SUM({N1895, N1894, N1893, N1892, N1891, N1890, 
        N1889, N1888, N1887, N1886}) );
  fpu_DW01_add_2 add_232 ( .A({1'b0, a_e}), .B({1'b0, b_e}), .CI(1'b0), .SUM({
        N936, N935, N934, N933, N932, N931, N930, N929, N928}) );
  fpu_DW01_inc_3 r392 ( .A(tmp_m1[22:1]), .SUM({N2316, N2315, N2314, N2313, 
        N2312, N2311, N2310, N2309, N2308, N2307, N2306, N2305, N2304, N2303, 
        N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295}) );
  fpu_DW01_inc_4 r391 ( .A(tmp_m1[23:2]), .SUM({N2264, N2263, N2262, N2261, 
        N2260, N2259, N2258, N2257, N2256, N2255, N2254, N2253, N2252, N2251, 
        N2250, N2249, N2248, N2247, N2246, N2245, N2244, N2243}) );
  fpu_DW01_inc_5 r390 ( .A(tmp_e1[7:0]), .SUM({N2242, N2241, N2240, N2239, 
        N2238, N2237, N2236, N2235}) );
  fpu_DW01_inc_6 r387 ( .A(tmp_m1), .SUM({N2450, N2228, N2227, N2226, N2225, 
        N2224, N2223, N2222, N2221, N2220, N2219, N2218, N2217, N2216, N2215, 
        N2214, N2213, N2212, N2211, N2210, N2209, N2208, N2207, N2206, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23}) );
  fpu_DW01_sub_24 r351 ( .A({1'b0, a_m[23], n1464, n1505, a_m[20], n1465, 
        n1506, n1472, n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, 
        a_m[9], n1480, n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0]}), .B({1'b0, n1467, b_m[22], n1938, b_m[20:18], n1936, n1934, b_m[15:14], 
        n1411, b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], n1930, b_m[1], 
        n1928}), .CI(1'b0), .DIFF({N483, N482, N481, N480, N479, N478, N477, 
        N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, 
        N464, N463, N462, N461, N460, N459}) );
  fpu_DW01_sub_25 r350 ( .A({1'b0, n1467, b_m[22], n1938, b_m[20:18], n1936, 
        n1934, b_m[15:14], n1410, b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], 
        n1930, b_m[1], n1928}), .B({1'b0, a_m[23], n1464, n1505, a_m[20], 
        n1465, n1506, n1472, n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, 
        a_m[9], n1480, n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0]}), .CI(1'b0), .DIFF({N458, N457, N456, N455, N454, N453, N452, N451, N450, 
        N449, N448, N447, N446, N445, N444, N443, N442, N441, N440, N439, N438, 
        N437, N436, N435, N434}) );
  fpu_DW01_sub_26 r349 ( .A({1'b0, a_m[23], n1464, n1505, a_m[20], n1465, 
        n1506, n1472, n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, 
        a_m[9], n1480, n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0]}), .B({1'b0, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, 
        N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, 
        N184}), .CI(1'b0), .DIFF({N432, N431, N430, N429, N428, N427, N426, 
        N425, N424, N423, N422, N421, N420, N419, N418, N417, N416, N415, N414, 
        N413, N412, N411, N410, N409, N408}) );
  fpu_DW01_sub_27 r348 ( .A({1'b0, n1467, b_m[22], n1938, b_m[20:18], n1936, 
        n1934, b_m[15:14], n1410, b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], 
        n1930, b_m[1], n1928}), .B({1'b0, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, 
        N131, N130, N129, N128, N127, N126}), .CI(1'b0), .DIFF({N374, N373, 
        N372, N371, N370, N369, N368, N367, N366, N365, N364, N363, N362, N361, 
        N360, N359, N358, N357, N356, N355, N354, N353, N352, N351, N350}) );
  fpu_DW01_add_3 r347 ( .A({1'b0, a_m[23], n1464, n1505, a_m[20], n1465, n1506, 
        n1472, n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, a_m[9], 
        n1480, n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0]}), .B({
        1'b0, n1467, b_m[22], n1938, b_m[20:18], n1936, n1934, b_m[15:14], 
        n1411, b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], n1930, b_m[1], 
        n1928}), .CI(1'b0), .SUM({N258, N257, N256, N255, N254, N253, N252, 
        N251, N250, N249, N248, N247, N246, N245, N244, N243, N242, N241, N240, 
        N239, N238, N237, N236, N235, N234}) );
  fpu_DW01_add_4 r346 ( .A({1'b0, a_m[23], n1464, n1505, a_m[20], n1465, n1506, 
        n1472, n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, a_m[9], 
        n1480, n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0]}), .B({
        1'b0, N207, N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, 
        N196, N195, N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, 
        N184}), .CI(1'b0), .SUM({N232, N231, N230, N229, N228, N227, N226, 
        N225, N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, 
        N213, N212, N211, N210, N209, N208}) );
  fpu_DW_rash_0 r345 ( .A({n1467, b_m[22], n1938, b_m[20:18], n1936, n1934, 
        b_m[15:14], n1410, b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], n1930, 
        b_m[1], n1928}), .DATA_TC(1'b0), .SH({N183, N182, N181, N180, N179, 
        N178, N177, N176}), .SH_TC(1'b0), .B({N207, N206, N205, N204, N203, 
        N202, N201, N200, N199, N198, N197, N196, N195, N194, N193, N192, N191, 
        N190, N189, N188, N187, N186, N185, N184}) );
  fpu_DW01_sub_28 r344 ( .A({1'b0, a_e}), .B({1'b0, b_e}), .CI(1'b0), .DIFF({
        N993, N183, N182, N181, N180, N179, N178, N177, N176}) );
  fpu_DW01_add_5 r343 ( .A({1'b0, n1467, b_m[22], n1938, b_m[20:18], n1936, 
        n1934, b_m[15:14], n1410, b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], 
        n1930, b_m[1], n1928}), .B({1'b0, N149, N148, N147, N146, N145, N144, 
        N143, N142, N141, N140, N139, N138, N137, N136, N135, N134, N133, N132, 
        N131, N130, N129, N128, N127, N126}), .CI(1'b0), .SUM({N174, N173, 
        N172, N171, N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, 
        N160, N159, N158, N157, N156, N155, N154, N153, N152, N151, N150}) );
  fpu_DW_rash_1 r342 ( .A({a_m[23], n1464, n1505, a_m[20], n1465, n1506, n1472, 
        n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, a_m[9], n1480, 
        n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0]}), .DATA_TC(
        1'b0), .SH({N125, N124, N123, N122, N121, N120, N119, N118}), .SH_TC(
        1'b0), .B({N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, 
        N139, N138, N137, N136, N135, N134, N133, N132, N131, N130, N129, N128, 
        N127, N126}) );
  fpu_DW01_sub_29 r341 ( .A(b_e), .B(a_e), .CI(1'b0), .DIFF({N125, N124, N123, 
        N122, N121, N120, N119, N118}) );
  fpu_DW02_mult_0 mult_233 ( .A({a_m[23], n1464, n1505, a_m[20], n1465, n1506, 
        n1472, n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, a_m[9], 
        n1480, n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0]}), .B({
        n1467, b_m[22], n1938, b_m[20:18], n1936, n1934, b_m[15:14], n1411, 
        b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], n1930, b_m[1], n1928}), 
        .TC(1'b0), .PRODUCT({N984, N983, N982, N981, N980, N979, N978, N977, 
        N976, N975, N974, N973, N972, N971, N970, N969, N968, N967, N966, N965, 
        N964, N963, N962, N961, N960, N959, N958, N957, N956, N955, N954, N953, 
        N952, N951, N950, N949, N948, N947, N946, N945, N944, N943, N942, N941, 
        N940, N939, N938, N937}) );
  DFFARX1_RVT \b_m_reg[0]  ( .D(b[0]), .CLK(clk), .RSTB(n1975), .Q(b_m[0]) );
  fpu_DW_div_uns_2 div_243 ( .a({a_m[23], n1464, n1505, a_m[20], n1465, n1506, 
        n1472, n1488, n1460, n1507, n1489, n1508, a_m[11], n1481, a_m[9], 
        n1480, n1466, n1509, n1482, n1510, n1483, n1490, n1511, a_m[0], 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .b({
        n1467, b_m[22], n1938, b_m[20:18], n1936, n1934, b_m[15:14], n1409, 
        b_m[12:9], n1932, b_m[7:6], n1931, b_m[4:3], n1930, b_m[1], n1928}), 
        .quotient({N1040, N1039, N1038, N1037, N1036, N1035, N1034, N1033, 
        N1032, N1031, N1030, N1029, N1028, N1027, N1026, N1025, N1024, N1023, 
        N1022, N1021, N1020, N1019, N1018, N1017, N1016, N1015, N1014, N1013, 
        N1012, N1011, N1010, N1009, N1008, N1007, N1006, N1005, N1004, N1003, 
        N1002, N1001, N1000, N999, N998, N997, N996, N995, N994}) );
  DFFARX1_RVT \tmp_m0_reg[26]  ( .D(N1078), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[26]) );
  DFFARX1_RVT \tmp_m0_reg[25]  ( .D(n1441), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[25]), .QN(n1695) );
  DFFARX1_RVT \tmp_m0_reg[2]  ( .D(N1054), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[2]), .QN(n1778) );
  DFFARX1_RVT \tmp_m0_reg[27]  ( .D(N1079), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[27]), .QN(n1475) );
  DFFARX1_RVT \tmp_m0_reg[28]  ( .D(N1080), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[28]), .QN(n1694) );
  DFFARX1_RVT \tmp_m0_reg[44]  ( .D(N1096), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[44]), .QN(n1795) );
  DFFARX1_RVT \tmp_m0_reg[16]  ( .D(N1068), .CLK(clk), .RSTB(n1962), .Q(
        tmp_m0[16]), .QN(n1792) );
  DFFARX1_RVT \tmp_m0_reg[15]  ( .D(N1067), .CLK(clk), .RSTB(n1962), .Q(
        tmp_m0[15]), .QN(n1791) );
  DFFARX1_RVT \tmp_m0_reg[14]  ( .D(N1066), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[14]), .QN(n1790) );
  DFFARX1_RVT \tmp_m0_reg[13]  ( .D(N1065), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[13]), .QN(n1613) );
  DFFARX1_RVT \tmp_m0_reg[36]  ( .D(N1088), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[36]), .QN(n1789) );
  DFFARX1_RVT \tmp_m0_reg[35]  ( .D(N1087), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[35]), .QN(n1787) );
  DFFARX1_RVT \tmp_m1_reg[44]  ( .D(N2109), .CLK(clk), .RSTB(n1971), .Q(
        tmp_m1[44]) );
  DFFX1_RVT \tmp_b_m0_reg[14]  ( .D(n1365), .CLK(clk), .Q(n1243) );
  DFFX1_RVT \tmp_b_m0_reg[2]  ( .D(n1341), .CLK(clk), .Q(n1231) );
  DFFARX1_RVT \tmp_m1_reg[47]  ( .D(N2112), .CLK(clk), .RSTB(n1971), .Q(
        tmp_m1[47]) );
  DFFARX1_RVT \tmp_m1_reg[46]  ( .D(n1630), .CLK(clk), .RSTB(n1971), .Q(
        tmp_m1[46]) );
  DFFARX1_RVT \tmp_m1_reg[45]  ( .D(n1688), .CLK(clk), .RSTB(n1971), .Q(
        tmp_m1[45]) );
  DFFARX1_RVT \tmp_m1_reg[1]  ( .D(N2066), .CLK(clk), .RSTB(n1967), .Q(
        tmp_m1[1]) );
  DFFARX1_RVT \tmp_m1_reg[17]  ( .D(n1587), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[17]) );
  DFFARX1_RVT \tmp_m1_reg[11]  ( .D(n1596), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[11]) );
  DFFARX1_RVT \tmp_m1_reg[6]  ( .D(N2071), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[6]) );
  DFFARX1_RVT \tmp_m1_reg[20]  ( .D(N2085), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[20]) );
  DFFARX1_RVT \tmp_m1_reg[15]  ( .D(N2080), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[15]) );
  DFFARX1_RVT \tmp_m1_reg[4]  ( .D(N2069), .CLK(clk), .RSTB(n1967), .Q(
        tmp_m1[4]) );
  DFFARX1_RVT \tmp_m1_reg[22]  ( .D(N2087), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[22]) );
  DFFARX1_RVT \tmp_m1_reg[21]  ( .D(N2086), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[21]) );
  DFFARX1_RVT \tmp_m1_reg[16]  ( .D(N2081), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[16]) );
  DFFARX1_RVT \tmp_m1_reg[10]  ( .D(n1622), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[10]) );
  DFFARX1_RVT \tmp_m1_reg[5]  ( .D(n1744), .CLK(clk), .RSTB(n1967), .Q(
        tmp_m1[5]) );
  DFFARX1_RVT \tmp_m1_reg[18]  ( .D(n1589), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[18]) );
  DFFARX1_RVT \tmp_m1_reg[12]  ( .D(n1628), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[12]) );
  DFFARX1_RVT \tmp_m1_reg[7]  ( .D(N2072), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[7]) );
  DFFARX1_RVT \tmp_m1_reg[14]  ( .D(N2079), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[14]) );
  DFFARX1_RVT \tmp_m1_reg[9]  ( .D(N2074), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[9]) );
  DFFARX1_RVT \tmp_m1_reg[3]  ( .D(N2068), .CLK(clk), .RSTB(n1967), .Q(
        tmp_m1[3]) );
  DFFARX1_RVT \tmp_m1_reg[19]  ( .D(N2084), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[19]) );
  DFFARX1_RVT \tmp_m1_reg[13]  ( .D(N2078), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[13]) );
  DFFARX1_RVT \tmp_m1_reg[8]  ( .D(N2073), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[8]) );
  DFFARX1_RVT \tmp_m1_reg[24]  ( .D(N2089), .CLK(clk), .RSTB(n1967), .Q(
        tmp_m1[24]) );
  DFFARX1_RVT \tmp_m1_reg[43]  ( .D(N2108), .CLK(clk), .RSTB(n1971), .Q(
        tmp_m1[43]) );
  DFFARX1_RVT \tmp_m1_reg[42]  ( .D(N2107), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[42]) );
  DFFARX1_RVT \tmp_m1_reg[41]  ( .D(N2106), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[41]) );
  DFFARX1_RVT \tmp_m1_reg[40]  ( .D(N2105), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[40]) );
  DFFARX1_RVT \tmp_m1_reg[39]  ( .D(N2104), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[39]) );
  DFFARX1_RVT \tmp_m1_reg[38]  ( .D(N2103), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[38]) );
  DFFARX1_RVT \tmp_m1_reg[37]  ( .D(N2102), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[37]) );
  DFFARX1_RVT \tmp_m1_reg[36]  ( .D(N2101), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[36]) );
  DFFARX1_RVT \tmp_m1_reg[35]  ( .D(N2100), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[35]) );
  DFFARX1_RVT \tmp_m1_reg[34]  ( .D(N2099), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[34]) );
  DFFARX1_RVT \tmp_m1_reg[33]  ( .D(N2098), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[33]) );
  DFFARX1_RVT \tmp_m1_reg[32]  ( .D(n1704), .CLK(clk), .RSTB(n1970), .Q(
        tmp_m1[32]) );
  DFFARX1_RVT \tmp_m1_reg[31]  ( .D(N2096), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[31]) );
  DFFARX1_RVT \tmp_m1_reg[30]  ( .D(n1720), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[30]) );
  DFFARX1_RVT \tmp_m1_reg[29]  ( .D(N2094), .CLK(clk), .RSTB(n1969), .Q(
        tmp_m1[29]) );
  DFFARX1_RVT \tmp_m1_reg[28]  ( .D(N2093), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[28]) );
  DFFARX1_RVT \tmp_m1_reg[27]  ( .D(N2092), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[27]) );
  DFFARX1_RVT \tmp_m1_reg[26]  ( .D(N2091), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[26]) );
  DFFARX1_RVT \tmp_m1_reg[2]  ( .D(N2067), .CLK(clk), .RSTB(n1967), .Q(
        tmp_m1[2]) );
  DFFARX1_RVT \tmp_m1_reg[25]  ( .D(N2090), .CLK(clk), .RSTB(n1968), .Q(
        tmp_m1[25]) );
  DFFARX1_RVT \tmp_e1_reg[8]  ( .D(N2063), .CLK(clk), .RSTB(n1967), .Q(
        tmp_e1[8]) );
  DFFARX1_RVT \tmp_e1_reg[9]  ( .D(N2064), .CLK(clk), .RSTB(n1967), .Q(
        tmp_e1[9]), .QN(n1784) );
  DFFARX1_RVT \tmp_e1_reg[3]  ( .D(N2058), .CLK(clk), .RSTB(n1966), .Q(
        tmp_e1[3]), .QN(n1181) );
  DFFARX1_RVT \tmp_e1_reg[6]  ( .D(N2061), .CLK(clk), .RSTB(n1966), .Q(
        tmp_e1[6]), .QN(n1184) );
  DFFARX1_RVT \tmp_e1_reg[2]  ( .D(n1450), .CLK(clk), .RSTB(n1966), .Q(
        tmp_e1[2]), .QN(n1180) );
  DFFARX1_RVT \tmp_e1_reg[7]  ( .D(N2062), .CLK(clk), .RSTB(n1970), .Q(
        tmp_e1[7]), .QN(n1185) );
  DFFARX1_RVT \tmp_e1_reg[5]  ( .D(N2060), .CLK(clk), .RSTB(n1966), .Q(
        tmp_e1[5]), .QN(n1183) );
  DFFARX1_RVT \tmp_e1_reg[4]  ( .D(N2059), .CLK(clk), .RSTB(n1966), .Q(
        tmp_e1[4]), .QN(n1182) );
  DFFARX1_RVT \tmp_e1_reg[1]  ( .D(n1728), .CLK(clk), .RSTB(n1966), .Q(
        tmp_e1[1]), .QN(n1179) );
  DFFARX1_RVT \tmp_e1_reg[0]  ( .D(N2055), .CLK(clk), .RSTB(n1966), .Q(
        tmp_e1[0]), .QN(n1178) );
  DFFARX1_RVT a_s_reg ( .D(a[31]), .CLK(clk), .RSTB(n1973), .Q(n1605) );
  DFFARX1_RVT \sel_0_reg[1]  ( .D(sel[1]), .CLK(clk), .RSTB(n1962), .Q(
        sel_0[1]), .QN(n1516) );
  DFFARX1_RVT b_s_reg ( .D(b[31]), .CLK(clk), .RSTB(n1972), .Q(n1609), .QN(
        n1398) );
  DFFARX1_RVT \sel_1_reg[0]  ( .D(sel_0[0]), .CLK(clk), .RSTB(n1972), .Q(
        sel_1[0]) );
  DFFARX1_RVT \sel_1_reg[1]  ( .D(sel_0[1]), .CLK(clk), .RSTB(n1960), .Q(
        sel_1[1]), .QN(n1560) );
  DFFARX1_RVT \tmp_m0_reg[47]  ( .D(N1099), .CLK(clk), .RSTB(n1971), .Q(
        tmp_m0[47]), .QN(n1561) );
  DFFARX1_RVT \tmp_m0_reg[45]  ( .D(N1097), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[45]), .QN(n1625) );
  DFFARX1_RVT \tmp_m0_reg[46]  ( .D(N1098), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[46]), .QN(n1606) );
  DFFARX1_RVT \tmp_m0_reg[5]  ( .D(N1057), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[5]), .QN(n1485) );
  DFFARX1_RVT \tmp_m0_reg[43]  ( .D(N1095), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[43]), .QN(n1615) );
  DFFARX1_RVT \tmp_m0_reg[9]  ( .D(N1061), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[9]) );
  DFFARX1_RVT \tmp_m0_reg[17]  ( .D(N1069), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[17]), .QN(n1468) );
  DFFARX1_RVT \tmp_m0_reg[18]  ( .D(N1070), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[18]), .QN(n1484) );
  DFFARX1_RVT \a_m_reg[18]  ( .D(a[18]), .CLK(clk), .RSTB(n1965), .Q(n1506), 
        .QN(n1571) );
  DFFARX1_RVT \a_m_reg[19]  ( .D(a[19]), .CLK(clk), .RSTB(n1965), .Q(n1465), 
        .QN(n1567) );
  DFFARX1_RVT \a_m_reg[20]  ( .D(a[20]), .CLK(clk), .RSTB(n1965), .Q(a_m[20]), 
        .QN(n1512) );
  DFFARX1_RVT \a_m_reg[17]  ( .D(a[17]), .CLK(clk), .RSTB(n1965), .Q(n1472), 
        .QN(n1566) );
  DFFARX1_RVT \a_m_reg[21]  ( .D(a[21]), .CLK(clk), .RSTB(n1966), .Q(n1505), 
        .QN(n1568) );
  DFFARX1_RVT \a_m_reg[22]  ( .D(a[22]), .CLK(clk), .RSTB(n1966), .Q(n1464), 
        .QN(n1572) );
  DFFARX1_RVT \a_m_reg[23]  ( .D(1'b1), .CLK(clk), .RSTB(n1966), .Q(a_m[23]), 
        .QN(n1515) );
  DFFARX1_RVT \tmp_e0_reg[7]  ( .D(N1048), .CLK(clk), .RSTB(n1972), .Q(n1525), 
        .QN(n1548) );
  DFFARX1_RVT \tmp_e0_reg[6]  ( .D(N1047), .CLK(clk), .RSTB(n1972), .Q(n1527), 
        .QN(n1547) );
  DFFARX1_RVT \tmp_e0_reg[5]  ( .D(N1046), .CLK(clk), .RSTB(n1972), .Q(n1526), 
        .QN(n1546) );
  DFFARX1_RVT \tmp_e0_reg[9]  ( .D(N1050), .CLK(clk), .RSTB(n1972), .QN(n1595)
         );
  DFFARX1_RVT \tmp_e0_reg[4]  ( .D(N1045), .CLK(clk), .RSTB(n1972), .QN(n1592)
         );
  DFFARX1_RVT \tmp_e0_reg[2]  ( .D(N1043), .CLK(clk), .RSTB(n1971), .QN(n1610)
         );
  DFFARX1_RVT \tmp_e0_reg[8]  ( .D(N1049), .CLK(clk), .RSTB(n1972), .Q(n1528), 
        .QN(n1594) );
  DFFARX1_RVT \tmp_e0_reg[3]  ( .D(N1044), .CLK(clk), .RSTB(n1972), .QN(n1591)
         );
  DFFARX1_RVT \tmp_e0_reg[1]  ( .D(N1042), .CLK(clk), .RSTB(n1971), .Q(N1188), 
        .QN(n1608) );
  DFFARX1_RVT \tmp_m0_reg[4]  ( .D(n1440), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[4]), .QN(n1497) );
  DFFARX1_RVT \tmp_m0_reg[3]  ( .D(N1055), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[3]), .QN(n1478) );
  DFFARX1_RVT \tmp_m0_reg[1]  ( .D(n1452), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[1]), .QN(n1462) );
  DFFARX1_RVT \a_m_reg[12]  ( .D(a[12]), .CLK(clk), .RSTB(n1965), .Q(n1508), 
        .QN(n1575) );
  DFFARX1_RVT \a_m_reg[11]  ( .D(a[11]), .CLK(clk), .RSTB(n1965), .Q(a_m[11]), 
        .QN(n1514) );
  DFFARX1_RVT \b_e_reg[7]  ( .D(b[30]), .CLK(clk), .RSTB(n1973), .Q(b_e[7]) );
  DFFARX1_RVT \b_m_reg[2]  ( .D(b[2]), .CLK(clk), .RSTB(n1962), .QN(n1573) );
  DFFARX1_RVT \b_m_reg[5]  ( .D(b[5]), .CLK(clk), .RSTB(n1962), .QN(n1416) );
  DFFARX1_RVT \b_m_reg[6]  ( .D(b[6]), .CLK(clk), .RSTB(n1962), .Q(b_m[6]) );
  DFFARX1_RVT \b_m_reg[4]  ( .D(b[4]), .CLK(clk), .RSTB(n1962), .Q(b_m[4]) );
  DFFARX1_RVT \b_m_reg[1]  ( .D(b[1]), .CLK(clk), .RSTB(n1962), .Q(b_m[1]) );
  DFFARX1_RVT \b_m_reg[20]  ( .D(b[20]), .CLK(clk), .RSTB(n1963), .Q(b_m[20])
         );
  DFFARX1_RVT \b_m_reg[17]  ( .D(b[17]), .CLK(clk), .RSTB(n1963), .Q(b_m[17])
         );
  DFFARX1_RVT \b_m_reg[18]  ( .D(b[18]), .CLK(clk), .RSTB(n1963), .Q(b_m[18])
         );
  DFFARX1_RVT \b_m_reg[21]  ( .D(b[21]), .CLK(clk), .RSTB(n1964), .Q(b_m[21])
         );
  DFFARX1_RVT \b_m_reg[22]  ( .D(b[22]), .CLK(clk), .RSTB(n1964), .Q(b_m[22])
         );
  DFFARX1_RVT \b_m_reg[23]  ( .D(1'b1), .CLK(clk), .RSTB(n1964), .Q(n1467), 
        .QN(n1574) );
  DFFARX1_RVT \b_e_reg[5]  ( .D(b[28]), .CLK(clk), .RSTB(n1973), .Q(b_e[5]), 
        .QN(n1537) );
  DFFARX1_RVT \b_e_reg[3]  ( .D(b[26]), .CLK(clk), .RSTB(n1973), .Q(b_e[3]), 
        .QN(n1536) );
  DFFARX1_RVT \a_e_reg[4]  ( .D(a[27]), .CLK(clk), .RSTB(n1974), .Q(a_e[4]), 
        .QN(n1261) );
  DFFARX1_RVT \b_e_reg[4]  ( .D(b[27]), .CLK(clk), .RSTB(n1973), .Q(b_e[4]) );
  DFFARX1_RVT \b_e_reg[6]  ( .D(b[29]), .CLK(clk), .RSTB(n1973), .Q(b_e[6]), 
        .QN(n1535) );
  DFFARX1_RVT \a_m_reg[2]  ( .D(a[2]), .CLK(clk), .RSTB(n1964), .Q(n1490), 
        .QN(n1581) );
  DFFARX1_RVT \a_m_reg[5]  ( .D(a[5]), .CLK(clk), .RSTB(n1964), .Q(n1482), 
        .QN(n1563) );
  DFFARX1_RVT \a_m_reg[6]  ( .D(a[6]), .CLK(clk), .RSTB(n1964), .Q(n1509), 
        .QN(n1577) );
  DFFARX1_RVT \a_m_reg[3]  ( .D(a[3]), .CLK(clk), .RSTB(n1964), .Q(n1483), 
        .QN(n1562) );
  DFFARX1_RVT \a_m_reg[4]  ( .D(a[4]), .CLK(clk), .RSTB(n1964), .Q(n1510), 
        .QN(n1576) );
  DFFARX1_RVT \a_m_reg[0]  ( .D(a[0]), .CLK(clk), .RSTB(n1964), .Q(a_m[0]), 
        .QN(n1517) );
  DFFARX1_RVT \a_m_reg[1]  ( .D(a[1]), .CLK(clk), .RSTB(n1964), .Q(n1511), 
        .QN(n1582) );
  DFFARX1_RVT \a_e_reg[2]  ( .D(a[25]), .CLK(clk), .RSTB(n1973), .Q(a_e[2]), 
        .QN(n1257) );
  DFFARX1_RVT \b_e_reg[2]  ( .D(b[25]), .CLK(clk), .RSTB(n1973), .Q(b_e[2]) );
  DFFARX1_RVT \tmp_m0_reg[10]  ( .D(N1062), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[10]), .QN(n1469) );
  DFFARX1_RVT \b_m_reg[11]  ( .D(b[11]), .CLK(clk), .RSTB(n1963), .Q(b_m[11])
         );
  DFFARX1_RVT \tmp_m0_reg[6]  ( .D(N1058), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[6]), .QN(n1494) );
  DFFARX1_RVT \a_m_reg[14]  ( .D(a[14]), .CLK(clk), .RSTB(n1965), .Q(n1507), 
        .QN(n1570) );
  DFFARX1_RVT \a_m_reg[13]  ( .D(a[13]), .CLK(clk), .RSTB(n1965), .Q(n1489), 
        .QN(n1569) );
  DFFARX1_RVT \a_m_reg[15]  ( .D(a[15]), .CLK(clk), .RSTB(n1965), .Q(n1460), 
        .QN(n1565) );
  DFFARX1_RVT \a_m_reg[16]  ( .D(a[16]), .CLK(clk), .RSTB(n1965), .Q(n1488), 
        .QN(n1579) );
  DFFARX1_RVT \a_m_reg[10]  ( .D(a[10]), .CLK(clk), .RSTB(n1965), .Q(n1481), 
        .QN(n1580) );
  DFFARX1_RVT \a_m_reg[8]  ( .D(a[8]), .CLK(clk), .RSTB(n1964), .Q(n1480), 
        .QN(n1578) );
  DFFARX1_RVT \a_m_reg[9]  ( .D(a[9]), .CLK(clk), .RSTB(n1965), .Q(a_m[9]), 
        .QN(n1513) );
  DFFARX1_RVT \a_m_reg[7]  ( .D(a[7]), .CLK(clk), .RSTB(n1964), .Q(n1466), 
        .QN(n1564) );
  DFFARX1_RVT \b_m_reg[14]  ( .D(b[14]), .CLK(clk), .RSTB(n1963), .Q(b_m[14])
         );
  DFFARX1_RVT \b_m_reg[15]  ( .D(b[15]), .CLK(clk), .RSTB(n1963), .Q(b_m[15])
         );
  DFFARX1_RVT \b_m_reg[16]  ( .D(b[16]), .CLK(clk), .RSTB(n1963), .Q(b_m[16])
         );
  DFFARX1_RVT \tmp_m0_reg[42]  ( .D(N1094), .CLK(clk), .RSTB(n1958), .Q(
        tmp_m0[42]), .QN(n1611) );
  DFFARX1_RVT \b_m_reg[12]  ( .D(b[12]), .CLK(clk), .RSTB(n1963), .Q(b_m[12])
         );
  DFFARX1_RVT \b_m_reg[13]  ( .D(b[13]), .CLK(clk), .RSTB(n1963), .Q(b_m[13])
         );
  DFFARX1_RVT \tmp_m0_reg[11]  ( .D(N1063), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[11]) );
  DFFARX1_RVT \tmp_m0_reg[23]  ( .D(N1075), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[23]), .QN(n1585) );
  DFFARX1_RVT \tmp_m0_reg[22]  ( .D(N1074), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[22]), .QN(n1474) );
  DFFARX1_RVT \tmp_m0_reg[20]  ( .D(N1072), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[20]), .QN(n1518) );
  DFFARX1_RVT \tmp_m0_reg[19]  ( .D(N1071), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[19]), .QN(n1492) );
  DFFARX1_RVT \tmp_m0_reg[7]  ( .D(N1059), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[7]) );
  DFFARX1_RVT \tmp_m0_reg[8]  ( .D(n1443), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[8]) );
  DFFARX1_RVT \tmp_m0_reg[37]  ( .D(N1089), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[37]), .QN(n1496) );
  DFFARX1_RVT \tmp_m0_reg[41]  ( .D(N1093), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[41]), .QN(n1612) );
  DFFARX1_RVT \tmp_m0_reg[38]  ( .D(N1090), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[38]), .QN(n1520) );
  DFFARX1_RVT \tmp_m0_reg[40]  ( .D(N1092), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[40]), .QN(n1461) );
  DFFARX1_RVT \tmp_m0_reg[39]  ( .D(N1091), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[39]), .QN(n1476) );
  DFFARX1_RVT \tmp_m0_reg[33]  ( .D(N1085), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[33]), .QN(n1470) );
  DFFARX1_RVT \tmp_m0_reg[32]  ( .D(N1084), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[32]), .QN(n1486) );
  DFFARX1_RVT \tmp_m0_reg[34]  ( .D(N1086), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[34]), .QN(n1623) );
  DFFARX1_RVT \tmp_m0_reg[12]  ( .D(N1064), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[12]), .QN(n1473) );
  DFFARX1_RVT \tmp_m0_reg[31]  ( .D(N1083), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[31]), .QN(n1545) );
  DFFARX1_RVT \tmp_m0_reg[30]  ( .D(N1082), .CLK(clk), .RSTB(n1959), .Q(
        tmp_m0[30]), .QN(n1690) );
  DFFARX1_RVT \tmp_m0_reg[29]  ( .D(N1081), .CLK(clk), .RSTB(n1960), .Q(
        tmp_m0[29]), .QN(n1504) );
  DFFARX1_RVT \b_m_reg[10]  ( .D(b[10]), .CLK(clk), .RSTB(n1963), .Q(b_m[10])
         );
  DFFARX1_RVT \b_m_reg[9]  ( .D(b[9]), .CLK(clk), .RSTB(n1963), .Q(b_m[9]) );
  DFFARX1_RVT \b_m_reg[8]  ( .D(b[8]), .CLK(clk), .RSTB(n1962), .Q(b_m[8]) );
  DFFARX1_RVT \b_m_reg[7]  ( .D(b[7]), .CLK(clk), .RSTB(n1962), .Q(b_m[7]) );
  DFFARX1_RVT \b_e_reg[0]  ( .D(b[23]), .CLK(clk), .RSTB(n1972), .Q(b_e[0]), 
        .QN(n1539) );
  DFFARX1_RVT \b_e_reg[1]  ( .D(b[24]), .CLK(clk), .RSTB(n1972), .Q(b_e[1]), 
        .QN(n1538) );
  DFFARX1_RVT \y_reg[31]  ( .D(N2800), .CLK(clk), .RSTB(n1966), .Q(y[31]) );
  DFFARX1_RVT \y_reg[30]  ( .D(N2799), .CLK(clk), .RSTB(n1966), .Q(y[30]) );
  DFFARX1_RVT \y_reg[29]  ( .D(N2798), .CLK(clk), .RSTB(n1967), .Q(y[29]) );
  DFFARX1_RVT \y_reg[28]  ( .D(N2797), .CLK(clk), .RSTB(n1967), .Q(y[28]) );
  DFFARX1_RVT \y_reg[27]  ( .D(N2796), .CLK(clk), .RSTB(n1967), .Q(y[27]) );
  DFFARX1_RVT \y_reg[26]  ( .D(N2795), .CLK(clk), .RSTB(n1974), .Q(y[26]) );
  DFFARX1_RVT \y_reg[25]  ( .D(N2794), .CLK(clk), .RSTB(n1974), .Q(y[25]) );
  DFFARX1_RVT \y_reg[24]  ( .D(N2793), .CLK(clk), .RSTB(n1973), .Q(y[24]) );
  DFFARX1_RVT \y_reg[23]  ( .D(N2792), .CLK(clk), .RSTB(n1974), .Q(y[23]) );
  DFFARX1_RVT \y_reg[22]  ( .D(N2791), .CLK(clk), .RSTB(n1974), .Q(y[22]) );
  DFFARX1_RVT \y_reg[21]  ( .D(N2790), .CLK(clk), .RSTB(n1974), .Q(y[21]) );
  DFFARX1_RVT \y_reg[20]  ( .D(N2789), .CLK(clk), .RSTB(n1974), .Q(y[20]) );
  DFFARX1_RVT \y_reg[19]  ( .D(N2788), .CLK(clk), .RSTB(n1974), .Q(y[19]) );
  DFFARX1_RVT \y_reg[18]  ( .D(N2787), .CLK(clk), .RSTB(n1974), .Q(y[18]) );
  DFFARX1_RVT \y_reg[17]  ( .D(N2786), .CLK(clk), .RSTB(n1974), .Q(y[17]) );
  DFFARX1_RVT \y_reg[16]  ( .D(N2785), .CLK(clk), .RSTB(n1975), .Q(y[16]) );
  DFFARX1_RVT \y_reg[15]  ( .D(N2784), .CLK(clk), .RSTB(n1975), .Q(y[15]) );
  DFFARX1_RVT \y_reg[14]  ( .D(N2783), .CLK(clk), .RSTB(n1975), .Q(y[14]) );
  DFFARX1_RVT \y_reg[13]  ( .D(N2782), .CLK(clk), .RSTB(n1974), .Q(y[13]) );
  DFFARX1_RVT \y_reg[12]  ( .D(N2781), .CLK(clk), .RSTB(n1961), .Q(y[12]) );
  DFFARX1_RVT \y_reg[11]  ( .D(N2780), .CLK(clk), .RSTB(n1957), .Q(y[11]) );
  DFFARX1_RVT \y_reg[10]  ( .D(N2779), .CLK(clk), .RSTB(n1957), .Q(y[10]) );
  DFFARX1_RVT \y_reg[9]  ( .D(N2778), .CLK(clk), .RSTB(n1957), .Q(y[9]) );
  DFFARX1_RVT \y_reg[8]  ( .D(N2777), .CLK(clk), .RSTB(n1957), .Q(y[8]) );
  DFFARX1_RVT \y_reg[7]  ( .D(N2776), .CLK(clk), .RSTB(n1957), .Q(y[7]) );
  DFFARX1_RVT \y_reg[6]  ( .D(N2775), .CLK(clk), .RSTB(n1957), .Q(y[6]) );
  DFFARX1_RVT \y_reg[5]  ( .D(N2774), .CLK(clk), .RSTB(n1957), .Q(y[5]) );
  DFFARX1_RVT \y_reg[4]  ( .D(N2773), .CLK(clk), .RSTB(n1957), .Q(y[4]) );
  DFFARX1_RVT \y_reg[3]  ( .D(N2772), .CLK(clk), .RSTB(n1957), .Q(y[3]) );
  DFFARX1_RVT \y_reg[2]  ( .D(N2771), .CLK(clk), .RSTB(n1957), .Q(y[2]) );
  DFFARX1_RVT \y_reg[1]  ( .D(N2770), .CLK(clk), .RSTB(n1957), .Q(y[1]) );
  DFFARX1_RVT \y_reg[0]  ( .D(N2769), .CLK(clk), .RSTB(n1958), .Q(y[0]) );
  DFFARX1_RVT tmp_s0_reg ( .D(N1051), .CLK(clk), .RSTB(n1971), .Q(tmp_s0) );
  DFFARX1_RVT err_reg ( .D(N2801), .CLK(clk), .RSTB(n1972), .Q(err) );
  DFFARX1_RVT overflow_reg ( .D(N2768), .CLK(clk), .RSTB(n1958), .Q(overflow)
         );
  DFFARX2_RVT \b_m_reg[19]  ( .D(b[19]), .CLK(clk), .RSTB(n1963), .Q(b_m[19])
         );
  DFFX1_RVT tmp_b_s0_reg ( .D(n1271), .CLK(clk), .Q(n1187) );
  DFFX1_RVT \tmp_a_e0_reg[7]  ( .D(n1397), .CLK(clk), .Q(n1266) );
  DFFX1_RVT \tmp_a_e0_reg[6]  ( .D(n1395), .CLK(clk), .Q(n1264) );
  DFFX1_RVT \tmp_a_e0_reg[5]  ( .D(n1393), .CLK(clk), .Q(n1262) );
  DFFX1_RVT \tmp_a_e0_reg[4]  ( .D(n1391), .CLK(clk), .Q(n1260) );
  DFFX1_RVT \tmp_a_e0_reg[3]  ( .D(n1389), .CLK(clk), .Q(n1258) );
  DFFX1_RVT tmp_a_s0_reg ( .D(n1335), .CLK(clk), .Q(n1227) );
  DFFX1_RVT \tmp_a_e0_reg[2]  ( .D(n1387), .CLK(clk), .Q(n1256) );
  DFFX1_RVT \tmp_a_e0_reg[1]  ( .D(n1385), .CLK(clk), .Q(n1254) );
  DFFX1_RVT \tmp_a_e0_reg[0]  ( .D(n1383), .CLK(clk), .Q(n1252) );
  DFFX1_RVT \tmp_b_e0_reg[7]  ( .D(n1287), .CLK(clk), .Q(n1202) );
  DFFX1_RVT \tmp_b_e0_reg[6]  ( .D(n1286), .CLK(clk), .Q(n1200) );
  DFFX1_RVT \tmp_b_e0_reg[5]  ( .D(n1285), .CLK(clk), .Q(n1198) );
  DFFX1_RVT \tmp_b_e0_reg[4]  ( .D(n1284), .CLK(clk), .Q(n1196) );
  DFFX1_RVT \tmp_b_e0_reg[3]  ( .D(n1283), .CLK(clk), .Q(n1194) );
  DFFX1_RVT \tmp_b_e0_reg[2]  ( .D(n1282), .CLK(clk), .Q(n1192) );
  DFFX1_RVT \tmp_b_e0_reg[1]  ( .D(n1281), .CLK(clk), .Q(n1190) );
  DFFX1_RVT \tmp_b_e0_reg[0]  ( .D(n1280), .CLK(clk), .Q(n1188) );
  DFFX1_RVT tmp_b_s1_reg ( .D(n1270), .CLK(clk), .Q(tmp_b_s1), .QN(n2471) );
  DFFX1_RVT tmp_a_s1_reg ( .D(n1334), .CLK(clk), .Q(tmp_a_s1), .QN(n2461) );
  DFFX1_RVT \tmp_b_m1_reg[2]  ( .D(n1340), .CLK(clk), .Q(tmp_b_m1[2]) );
  DFFX1_RVT \tmp_a_m1_reg[20]  ( .D(n1328), .CLK(clk), .Q(tmp_a_m1[20]) );
  DFFX1_RVT \tmp_a_m1_reg[13]  ( .D(n1314), .CLK(clk), .Q(tmp_a_m1[13]) );
  DFFX1_RVT \tmp_a_m1_reg[15]  ( .D(n1318), .CLK(clk), .Q(tmp_a_m1[15]) );
  DFFX1_RVT \tmp_a_m1_reg[18]  ( .D(n1324), .CLK(clk), .Q(tmp_a_m1[18]) );
  DFFX1_RVT \tmp_a_m1_reg[21]  ( .D(n1330), .CLK(clk), .Q(tmp_a_m1[21]) );
  DFFX1_RVT \tmp_a_m1_reg[12]  ( .D(n1312), .CLK(clk), .Q(tmp_a_m1[12]) );
  DFFX1_RVT \tmp_a_m1_reg[16]  ( .D(n1320), .CLK(clk), .Q(tmp_a_m1[16]) );
  DFFX1_RVT \tmp_a_m1_reg[0]  ( .D(n1288), .CLK(clk), .Q(tmp_a_m1[0]), .QN(
        n2463) );
  DFFX1_RVT \tmp_a_m1_reg[19]  ( .D(n1326), .CLK(clk), .Q(tmp_a_m1[19]) );
  DFFX1_RVT \tmp_a_m1_reg[9]  ( .D(n1306), .CLK(clk), .Q(tmp_a_m1[9]) );
  DFFX1_RVT \tmp_a_m1_reg[14]  ( .D(n1316), .CLK(clk), .Q(tmp_a_m1[14]) );
  DFFX1_RVT \tmp_a_m1_reg[5]  ( .D(n1298), .CLK(clk), .Q(tmp_a_m1[5]) );
  DFFX1_RVT \tmp_a_m1_reg[8]  ( .D(n1304), .CLK(clk), .Q(tmp_a_m1[8]) );
  DFFX1_RVT \tmp_b_m1_reg[5]  ( .D(n1346), .CLK(clk), .Q(tmp_b_m1[5]) );
  DFFX1_RVT \tmp_a_m1_reg[22]  ( .D(n1332), .CLK(clk), .Q(tmp_a_m1[22]) );
  DFFX1_RVT \tmp_a_m1_reg[17]  ( .D(n1322), .CLK(clk), .Q(tmp_a_m1[17]) );
  DFFX1_RVT \tmp_a_m1_reg[6]  ( .D(n1300), .CLK(clk), .Q(tmp_a_m1[6]) );
  DFFX1_RVT \tmp_a_m1_reg[2]  ( .D(n1292), .CLK(clk), .Q(tmp_a_m1[2]) );
  DFFX1_RVT \tmp_b_m1_reg[6]  ( .D(n1348), .CLK(clk), .Q(tmp_b_m1[6]) );
  DFFX1_RVT \tmp_a_m1_reg[4]  ( .D(n1296), .CLK(clk), .Q(tmp_a_m1[4]) );
  DFFX1_RVT \tmp_a_m1_reg[11]  ( .D(n1310), .CLK(clk), .Q(tmp_a_m1[11]) );
  DFFX1_RVT \tmp_a_m1_reg[3]  ( .D(n1294), .CLK(clk), .Q(tmp_a_m1[3]) );
  DFFX1_RVT \tmp_b_m1_reg[4]  ( .D(n1344), .CLK(clk), .Q(tmp_b_m1[4]) );
  DFFX1_RVT \tmp_b_m1_reg[20]  ( .D(n1376), .CLK(clk), .Q(tmp_b_m1[20]) );
  DFFX1_RVT \tmp_b_m1_reg[3]  ( .D(n1342), .CLK(clk), .Q(tmp_b_m1[3]) );
  DFFX1_RVT \tmp_a_e1_reg[6]  ( .D(n1394), .CLK(clk), .Q(tmp_a_e1[6]), .QN(
        n2451) );
  DFFX1_RVT \tmp_b_m1_reg[15]  ( .D(n1366), .CLK(clk), .Q(tmp_b_m1[15]) );
  DFFX1_RVT \tmp_a_m1_reg[7]  ( .D(n1302), .CLK(clk), .Q(tmp_a_m1[7]) );
  DFFX1_RVT \tmp_b_m1_reg[18]  ( .D(n1372), .CLK(clk), .Q(tmp_b_m1[18]) );
  DFFX1_RVT \tmp_b_m1_reg[8]  ( .D(n1352), .CLK(clk), .Q(tmp_b_m1[8]) );
  DFFX1_RVT \tmp_a_e1_reg[5]  ( .D(n1392), .CLK(clk), .Q(tmp_a_e1[5]), .QN(
        n2452) );
  DFFX1_RVT \tmp_a_e1_reg[4]  ( .D(n1390), .CLK(clk), .Q(tmp_a_e1[4]), .QN(
        n2453) );
  DFFX1_RVT \tmp_b_m1_reg[21]  ( .D(n1378), .CLK(clk), .Q(tmp_b_m1[21]) );
  DFFX1_RVT \tmp_b_m1_reg[12]  ( .D(n1360), .CLK(clk), .Q(tmp_b_m1[12]) );
  DFFX1_RVT \tmp_b_m1_reg[16]  ( .D(n1368), .CLK(clk), .Q(tmp_b_m1[16]) );
  DFFX1_RVT \tmp_b_m1_reg[19]  ( .D(n1374), .CLK(clk), .Q(tmp_b_m1[19]) );
  DFFX1_RVT \tmp_b_m1_reg[9]  ( .D(n1354), .CLK(clk), .Q(tmp_b_m1[9]) );
  DFFX1_RVT \tmp_b_m1_reg[13]  ( .D(n1362), .CLK(clk), .Q(tmp_b_m1[13]) );
  DFFX1_RVT \tmp_b_m1_reg[1]  ( .D(n1338), .CLK(clk), .Q(tmp_b_m1[1]), .QN(
        n2420) );
  DFFX1_RVT \tmp_b_m1_reg[14]  ( .D(n1364), .CLK(clk), .Q(tmp_b_m1[14]) );
  DFFX1_RVT \tmp_a_e1_reg[3]  ( .D(n1388), .CLK(clk), .Q(tmp_a_e1[3]), .QN(
        n2454) );
  DFFX1_RVT \tmp_a_m1_reg[10]  ( .D(n1308), .CLK(clk), .Q(tmp_a_m1[10]), .QN(
        n2462) );
  DFFX1_RVT \tmp_b_m1_reg[22]  ( .D(n1380), .CLK(clk), .Q(tmp_b_m1[22]) );
  DFFX1_RVT \tmp_b_m1_reg[17]  ( .D(n1370), .CLK(clk), .Q(tmp_b_m1[17]) );
  DFFX1_RVT \tmp_b_m1_reg[7]  ( .D(n1350), .CLK(clk), .Q(tmp_b_m1[7]) );
  DFFX1_RVT \tmp_a_e1_reg[7]  ( .D(n1396), .CLK(clk), .Q(tmp_a_e1[7]), .QN(
        n2446) );
  DFFX1_RVT \tmp_b_m1_reg[11]  ( .D(n1358), .CLK(clk), .Q(tmp_b_m1[11]) );
  DFFX1_RVT \tmp_b_m1_reg[10]  ( .D(n1356), .CLK(clk), .Q(tmp_b_m1[10]), .QN(
        n2459) );
  DFFX1_RVT \tmp_a_m1_reg[1]  ( .D(n1290), .CLK(clk), .Q(tmp_a_m1[1]), .QN(
        n2419) );
  DFFX1_RVT \tmp_b_e1_reg[6]  ( .D(n1278), .CLK(clk), .Q(tmp_b_e1[6]), .QN(
        n2466) );
  DFFX1_RVT \tmp_b_e1_reg[5]  ( .D(n1277), .CLK(clk), .Q(tmp_b_e1[5]), .QN(
        n2467) );
  DFFX1_RVT \tmp_b_e1_reg[4]  ( .D(n1276), .CLK(clk), .Q(tmp_b_e1[4]), .QN(
        n2468) );
  DFFX1_RVT \tmp_b_m1_reg[0]  ( .D(n1336), .CLK(clk), .Q(tmp_b_m1[0]), .QN(
        n2460) );
  DFFX1_RVT \tmp_b_e1_reg[0]  ( .D(n1272), .CLK(clk), .Q(tmp_b_e1[0]), .QN(
        n2384) );
  DFFX1_RVT \tmp_b_e1_reg[7]  ( .D(n1279), .CLK(clk), .Q(tmp_b_e1[7]), .QN(
        n2464) );
  DFFX1_RVT \tmp_b_e1_reg[3]  ( .D(n1275), .CLK(clk), .Q(tmp_b_e1[3]), .QN(
        n2469) );
  DFFX1_RVT \tmp_a_e1_reg[2]  ( .D(n1386), .CLK(clk), .Q(tmp_a_e1[2]), .QN(
        n2455) );
  DFFX1_RVT \tmp_b_e1_reg[2]  ( .D(n1274), .CLK(clk), .Q(tmp_b_e1[2]), .QN(
        n2470) );
  DFFX1_RVT \tmp_b_e1_reg[1]  ( .D(n1273), .CLK(clk), .Q(tmp_b_e1[1]), .QN(
        n2385) );
  DFFX1_RVT \tmp_a_e1_reg[0]  ( .D(n1382), .CLK(clk), .Q(tmp_a_e1[0]), .QN(
        n2457) );
  DFFX1_RVT \tmp_a_e1_reg[1]  ( .D(n1384), .CLK(clk), .Q(tmp_a_e1[1]), .QN(
        n2456) );
  DFFX1_RVT \sel_2_reg[1]  ( .D(n1269), .CLK(clk), .Q(\sel_2[1] ), .QN(n2474)
         );
  DFFX1_RVT \sel_2_reg[0]  ( .D(n1268), .CLK(clk), .Q(n1186), .QN(n2476) );
  DFFX1_RVT \tmp_b_m0_reg[12]  ( .D(n1361), .CLK(clk), .Q(n1241) );
  DFFX1_RVT \tmp_b_m0_reg[13]  ( .D(n1363), .CLK(clk), .Q(n1242) );
  DFFX1_RVT \tmp_b_m0_reg[11]  ( .D(n1359), .CLK(clk), .Q(n1240) );
  DFFX1_RVT \tmp_b_m0_reg[10]  ( .D(n1357), .CLK(clk), .Q(n1239) );
  DFFX1_RVT \tmp_b_m0_reg[0]  ( .D(n1337), .CLK(clk), .Q(n1229) );
  DFFX1_RVT \tmp_b_m0_reg[1]  ( .D(n1339), .CLK(clk), .Q(n1230) );
  DFFX1_RVT \tmp_b_m0_reg[22]  ( .D(n1381), .CLK(clk), .Q(n1251) );
  DFFX1_RVT \tmp_b_m0_reg[19]  ( .D(n1375), .CLK(clk), .Q(n1248) );
  DFFX1_RVT \tmp_a_m0_reg[20]  ( .D(n1329), .CLK(clk), .Q(n1224) );
  DFFX1_RVT \tmp_b_m0_reg[6]  ( .D(n1349), .CLK(clk), .Q(n1235) );
  DFFX1_RVT \tmp_b_m0_reg[4]  ( .D(n1345), .CLK(clk), .Q(n1233) );
  DFFX1_RVT \tmp_b_m0_reg[9]  ( .D(n1355), .CLK(clk), .Q(n1238) );
  DFFX1_RVT \tmp_b_m0_reg[7]  ( .D(n1351), .CLK(clk), .Q(n1236) );
  DFFX1_RVT \tmp_b_m0_reg[8]  ( .D(n1353), .CLK(clk), .Q(n1237) );
  DFFX1_RVT \tmp_b_m0_reg[3]  ( .D(n1343), .CLK(clk), .Q(n1232) );
  DFFX1_RVT \tmp_a_m0_reg[0]  ( .D(n1289), .CLK(clk), .Q(n1204) );
  DFFX1_RVT \tmp_a_m0_reg[14]  ( .D(n1317), .CLK(clk), .Q(n1218) );
  DFFX1_RVT \tmp_a_m0_reg[6]  ( .D(n1301), .CLK(clk), .Q(n1210) );
  DFFX1_RVT \tmp_a_m0_reg[5]  ( .D(n1299), .CLK(clk), .Q(n1209) );
  DFFX1_RVT \tmp_a_m0_reg[2]  ( .D(n1293), .CLK(clk), .Q(n1206) );
  DFFX1_RVT \tmp_b_m0_reg[21]  ( .D(n1379), .CLK(clk), .Q(n1250) );
  DFFX1_RVT \tmp_a_m0_reg[3]  ( .D(n1295), .CLK(clk), .Q(n1207) );
  DFFX1_RVT \tmp_b_m0_reg[20]  ( .D(n1377), .CLK(clk), .Q(n1249) );
  DFFX1_RVT \tmp_a_m0_reg[22]  ( .D(n1333), .CLK(clk), .Q(n1226) );
  DFFX1_RVT \tmp_a_m0_reg[18]  ( .D(n1325), .CLK(clk), .Q(n1222) );
  DFFX1_RVT \tmp_a_m0_reg[16]  ( .D(n1321), .CLK(clk), .Q(n1220) );
  DFFX1_RVT \tmp_a_m0_reg[4]  ( .D(n1297), .CLK(clk), .Q(n1208) );
  DFFX1_RVT \tmp_a_m0_reg[19]  ( .D(n1327), .CLK(clk), .Q(n1223) );
  DFFX1_RVT \tmp_a_m0_reg[17]  ( .D(n1323), .CLK(clk), .Q(n1221) );
  DFFX1_RVT \tmp_a_m0_reg[15]  ( .D(n1319), .CLK(clk), .Q(n1219) );
  DFFX1_RVT \tmp_a_m0_reg[9]  ( .D(n1307), .CLK(clk), .Q(n1213) );
  DFFX1_RVT \tmp_a_m0_reg[7]  ( .D(n1303), .CLK(clk), .Q(n1211) );
  DFFX1_RVT \tmp_a_m0_reg[8]  ( .D(n1305), .CLK(clk), .Q(n1212) );
  DFFX1_RVT \tmp_a_m0_reg[21]  ( .D(n1331), .CLK(clk), .Q(n1225) );
  DFFX1_RVT \tmp_b_m0_reg[5]  ( .D(n1347), .CLK(clk), .Q(n1234) );
  DFFX1_RVT \tmp_b_m0_reg[17]  ( .D(n1371), .CLK(clk), .Q(n1246) );
  DFFX1_RVT \tmp_b_m0_reg[15]  ( .D(n1367), .CLK(clk), .Q(n1244) );
  DFFX1_RVT \tmp_b_m0_reg[18]  ( .D(n1373), .CLK(clk), .Q(n1247) );
  DFFX1_RVT \tmp_b_m0_reg[16]  ( .D(n1369), .CLK(clk), .Q(n1245) );
  DFFX1_RVT \tmp_a_m0_reg[1]  ( .D(n1291), .CLK(clk), .Q(n1205) );
  DFFX1_RVT \tmp_a_m0_reg[12]  ( .D(n1313), .CLK(clk), .Q(n1216) );
  DFFX1_RVT \tmp_a_m0_reg[13]  ( .D(n1315), .CLK(clk), .Q(n1217) );
  DFFX1_RVT \tmp_a_m0_reg[11]  ( .D(n1311), .CLK(clk), .Q(n1215) );
  DFFX1_RVT \tmp_a_m0_reg[10]  ( .D(n1309), .CLK(clk), .Q(n1214) );
  DFFARX1_RVT tmp_s1_reg ( .D(tmp_s0), .CLK(clk), .RSTB(n1956), .QN(n2477) );
  DFFARX1_RVT \a_e_reg[7]  ( .D(a[30]), .CLK(clk), .RSTB(n1957), .Q(a_e[7]), 
        .QN(n1267) );
  DFFARX1_RVT \a_e_reg[6]  ( .D(a[29]), .CLK(clk), .RSTB(n1971), .Q(a_e[6]), 
        .QN(n1265) );
  DFFARX1_RVT \a_e_reg[1]  ( .D(a[24]), .CLK(clk), .RSTB(n1973), .Q(a_e[1]), 
        .QN(n1255) );
  DFFARX1_RVT \tmp_m0_reg[24]  ( .D(N1076), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[24]), .QN(n1559) );
  DFFARX1_RVT \a_e_reg[5]  ( .D(a[28]), .CLK(clk), .RSTB(n1974), .Q(a_e[5]) );
  DFFARX1_RVT \a_e_reg[3]  ( .D(a[26]), .CLK(clk), .RSTB(n1973), .Q(a_e[3]) );
  DFFARX1_RVT \a_e_reg[0]  ( .D(a[23]), .CLK(clk), .RSTB(n1973), .Q(a_e[0]) );
  DFFARX1_RVT \tmp_m0_reg[0]  ( .D(n1459), .CLK(clk), .RSTB(n1967), .Q(
        tmp_m0[0]), .QN(n1533) );
  DFFARX2_RVT \b_m_reg[3]  ( .D(b[3]), .CLK(clk), .RSTB(n1962), .Q(b_m[3]) );
  DFFARX1_RVT \sel_0_reg[0]  ( .D(sel[0]), .CLK(clk), .RSTB(n1962), .Q(
        sel_0[0]) );
  DFFARX1_RVT \tmp_e0_reg[0]  ( .D(N1041), .CLK(clk), .RSTB(n1955), .Q(N1129)
         );
  DFFARX1_RVT \tmp_m0_reg[21]  ( .D(N1073), .CLK(clk), .RSTB(n1961), .Q(
        tmp_m0[21]), .QN(n1493) );
  INVX4_RVT U1330 ( .A(n1405), .Y(n1402) );
  IBUFFX4_RVT U1331 ( .A(n1402), .Y(n1403) );
  IBUFFX32_RVT U1332 ( .A(n1404), .Y(n1405) );
  INVX2_RVT U1333 ( .A(n1458), .Y(n1404) );
  IBUFFX16_RVT U1334 ( .A(N1052), .Y(n1458) );
  INVX2_RVT U1335 ( .A(n1403), .Y(n1406) );
  IBUFFX4_RVT U1336 ( .A(n1406), .Y(n1407) );
  IBUFFX32_RVT U1337 ( .A(n1407), .Y(n1459) );
  IBUFFX4_RVT U1338 ( .A(b_m[13]), .Y(n1408) );
  INVX2_RVT U1339 ( .A(n1408), .Y(n1409) );
  INVX0_RVT U1340 ( .A(n1408), .Y(n1410) );
  INVX0_RVT U1341 ( .A(n1408), .Y(n1411) );
  INVX4_RVT U1342 ( .A(N2057), .Y(n1449) );
  INVX4_RVT U1343 ( .A(N2097), .Y(n1703) );
  IBUFFX16_RVT U1344 ( .A(n1686), .Y(n1728) );
  INVX4_RVT U1345 ( .A(n1685), .Y(n1686) );
  INVX1_RVT U1346 ( .A(n1933), .Y(n1932) );
  INVX1_RVT U1347 ( .A(n1912), .Y(n1911) );
  INVX1_RVT U1348 ( .A(n1424), .Y(n1896) );
  INVX1_RVT U1349 ( .A(n1891), .Y(n1897) );
  INVX1_RVT U1350 ( .A(n1424), .Y(n1901) );
  INVX1_RVT U1351 ( .A(n581), .Y(n1700) );
  INVX1_RVT U1352 ( .A(n1786), .Y(n1809) );
  INVX1_RVT U1353 ( .A(N1129), .Y(n1430) );
  INVX1_RVT U1354 ( .A(n967), .Y(n1759) );
  AO222X1_RVT U1355 ( .A1(N1745), .A2(n1862), .A3(N1321), .A4(n1812), .A5(
        n1610), .A6(n1895), .Y(n967) );
  INVX2_RVT U1356 ( .A(n1702), .Y(n1439) );
  NOR2X1_RVT U1357 ( .A1(n1002), .A2(n994), .Y(n870) );
  INVX1_RVT U1358 ( .A(n461), .Y(n2482) );
  AND4X1_RVT U1359 ( .A1(n543), .A2(n544), .A3(n542), .A4(n2129), .Y(n2130) );
  INVX0_RVT U1360 ( .A(n1809), .Y(n1811) );
  INVX1_RVT U1361 ( .A(n515), .Y(n1785) );
  INVX1_RVT U1362 ( .A(n501), .Y(n1804) );
  INVX1_RVT U1363 ( .A(n1767), .Y(n501) );
  AND2X1_RVT U1364 ( .A1(n2087), .A2(n2322), .Y(n1767) );
  INVX1_RVT U1365 ( .A(n2295), .Y(n2087) );
  NAND2X0_RVT U1366 ( .A1(n2099), .A2(n1484), .Y(n1495) );
  INVX1_RVT U1367 ( .A(n1543), .Y(n1793) );
  NAND2X0_RVT U1368 ( .A1(tmp_m0[15]), .A2(n1842), .Y(n402) );
  INVX1_RVT U1369 ( .A(n2293), .Y(n2095) );
  INVX1_RVT U1370 ( .A(n1150), .Y(n2438) );
  INVX1_RVT U1371 ( .A(n1176), .Y(n2324) );
  INVX1_RVT U1372 ( .A(n2367), .Y(n2371) );
  INVX1_RVT U1373 ( .A(n1698), .Y(n1699) );
  INVX1_RVT U1374 ( .A(n2091), .Y(n1698) );
  INVX1_RVT U1375 ( .A(n2078), .Y(n2091) );
  INVX1_RVT U1376 ( .A(n2089), .Y(n2088) );
  INVX1_RVT U1377 ( .A(n1419), .Y(n1641) );
  INVX1_RVT U1378 ( .A(n1423), .Y(n1639) );
  INVX1_RVT U1379 ( .A(n1422), .Y(n1637) );
  INVX1_RVT U1380 ( .A(n1421), .Y(n1635) );
  INVX1_RVT U1381 ( .A(n1420), .Y(n1633) );
  INVX1_RVT U1382 ( .A(n1418), .Y(n1643) );
  INVX1_RVT U1383 ( .A(n1417), .Y(n1645) );
  IBUFFX16_RVT U1384 ( .A(n534), .Y(n1715) );
  NAND4X0_RVT U1385 ( .A1(n536), .A2(n537), .A3(n538), .A4(n539), .Y(n534) );
  NAND4X0_RVT U1386 ( .A1(n525), .A2(n526), .A3(n527), .A4(n528), .Y(n523) );
  IBUFFX16_RVT U1387 ( .A(n509), .Y(n1730) );
  NAND4X0_RVT U1388 ( .A1(n511), .A2(n512), .A3(n513), .A4(n514), .Y(n509) );
  NAND2X0_RVT U1389 ( .A1(n1807), .A2(n1543), .Y(n576) );
  INVX1_RVT U1390 ( .A(n2294), .Y(n2108) );
  INVX1_RVT U1391 ( .A(n1424), .Y(n1900) );
  INVX1_RVT U1392 ( .A(n647), .Y(n2099) );
  INVX1_RVT U1393 ( .A(n1588), .Y(n1424) );
  INVX1_RVT U1394 ( .A(n1769), .Y(n1884) );
  INVX1_RVT U1395 ( .A(n1785), .Y(n1786) );
  INVX1_RVT U1396 ( .A(n426), .Y(n2113) );
  INVX1_RVT U1397 ( .A(n428), .Y(n2114) );
  INVX1_RVT U1398 ( .A(n1817), .Y(n1818) );
  NBUFFX2_RVT U1399 ( .A(n2296), .Y(n1813) );
  INVX1_RVT U1400 ( .A(n1898), .Y(n1892) );
  INVX1_RVT U1401 ( .A(n1807), .Y(n1808) );
  INVX1_RVT U1402 ( .A(n1424), .Y(n1898) );
  INVX1_RVT U1403 ( .A(n994), .Y(n2322) );
  MUX21X1_RVT U1404 ( .A1(n2017), .A2(n1144), .S0(sel_0[0]), .Y(n2018) );
  AO221X1_RVT U1405 ( .A1(N236), .A2(net32932), .A3(N210), .A4(net32938), .A5(
        n2115), .Y(n2116) );
  INVX1_RVT U1406 ( .A(n1540), .Y(n1862) );
  XNOR2X1_RVT U1407 ( .A1(n1605), .A2(n1398), .Y(n1147) );
  INVX1_RVT U1408 ( .A(n2106), .Y(n1447) );
  AO222X1_RVT U1409 ( .A1(N439), .A2(net32946), .A3(N355), .A4(net32952), .A5(
        N413), .A6(net27438), .Y(n2106) );
  INVX1_RVT U1410 ( .A(N1129), .Y(n1429) );
  NOR2X1_RVT U1411 ( .A1(n1584), .A2(n1853), .Y(n1433) );
  AO221X1_RVT U1412 ( .A1(n1608), .A2(n1864), .A3(N2036), .A4(n2317), .A5(n970), .Y(N2056) );
  OR2X1_RVT U1413 ( .A1(n1642), .A2(n1650), .Y(n932) );
  INVX1_RVT U1414 ( .A(n1641), .Y(n1642) );
  OR2X1_RVT U1415 ( .A1(n1640), .A2(n1652), .Y(n919) );
  INVX1_RVT U1416 ( .A(n1639), .Y(n1640) );
  OR2X1_RVT U1417 ( .A1(n1638), .A2(n1656), .Y(n893) );
  INVX1_RVT U1418 ( .A(n1637), .Y(n1638) );
  INVX1_RVT U1419 ( .A(n1608), .Y(n1909) );
  OR2X1_RVT U1420 ( .A1(n1636), .A2(n1654), .Y(n906) );
  INVX1_RVT U1421 ( .A(n1635), .Y(n1636) );
  OR2X1_RVT U1422 ( .A1(n1634), .A2(n1648), .Y(n945) );
  INVX1_RVT U1423 ( .A(n1633), .Y(n1634) );
  OR2X1_RVT U1424 ( .A1(n1644), .A2(n1660), .Y(n851) );
  INVX1_RVT U1425 ( .A(n1643), .Y(n1644) );
  OR2X1_RVT U1426 ( .A1(n1646), .A2(n1658), .Y(n880) );
  INVX1_RVT U1427 ( .A(n1645), .Y(n1646) );
  NBUFFX2_RVT U1428 ( .A(n2132), .Y(n1816) );
  INVX1_RVT U1429 ( .A(tmp_m0[28]), .Y(n2316) );
  OA222X1_RVT U1430 ( .A1(n1790), .A2(n1559), .A3(n580), .A4(n1497), .A5(n1892), .A6(n1803), .Y(n2196) );
  NAND2X0_RVT U1431 ( .A1(tmp_m0[8]), .A2(n2322), .Y(n1692) );
  INVX1_RVT U1432 ( .A(tmp_m0[8]), .Y(n2301) );
  INVX4_RVT U1433 ( .A(n2246), .Y(n1681) );
  OAI221X1_RVT U1434 ( .A1(n1786), .A2(n2291), .A3(n648), .A4(n2245), .A5(
        n2244), .Y(n1682) );
  INVX1_RVT U1435 ( .A(n1779), .Y(n1867) );
  INVX4_RVT U1436 ( .A(n2178), .Y(n1677) );
  INVX1_RVT U1437 ( .A(n1862), .Y(n1860) );
  INVX1_RVT U1438 ( .A(n1424), .Y(n1899) );
  OAI221X1_RVT U1439 ( .A1(n1691), .A2(n1485), .A3(n648), .A4(n2266), .A5(
        n2265), .Y(n1666) );
  NAND2X0_RVT U1440 ( .A1(tmp_m0[8]), .A2(n2322), .Y(n1691) );
  INVX4_RVT U1441 ( .A(n2269), .Y(n1665) );
  INVX1_RVT U1442 ( .A(n1878), .Y(n1877) );
  INVX4_RVT U1443 ( .A(n2182), .Y(n1673) );
  NBUFFX2_RVT U1444 ( .A(n2300), .Y(n1801) );
  INVX1_RVT U1445 ( .A(n1871), .Y(n1868) );
  INVX1_RVT U1446 ( .A(n1883), .Y(n1879) );
  OAI222X1_RVT U1447 ( .A1(n1806), .A2(n1462), .A3(n648), .A4(n2236), .A5(n515), .A6(n2287), .Y(n1670) );
  INVX4_RVT U1448 ( .A(n2237), .Y(n1669) );
  AOI221X1_RVT U1449 ( .A1(n2320), .A2(n488), .A3(tmp_m0[42]), .A4(n1863), 
        .A5(n489), .Y(n484) );
  INVX1_RVT U1450 ( .A(n1752), .Y(n1631) );
  INVX1_RVT U1451 ( .A(n1753), .Y(n1752) );
  INVX1_RVT U1452 ( .A(n1435), .Y(n1753) );
  INVX1_RVT U1453 ( .A(n1890), .Y(n1885) );
  INVX1_RVT U1454 ( .A(n2322), .Y(n1794) );
  NOR2X1_RVT U1455 ( .A1(n1853), .A2(n1739), .Y(n1741) );
  INVX1_RVT U1456 ( .A(n495), .Y(n1739) );
  INVX1_RVT U1457 ( .A(n2116), .Y(n1455) );
  INVX1_RVT U1458 ( .A(n2288), .Y(n2315) );
  NAND3X0_RVT U1459 ( .A1(n1593), .A2(n2123), .A3(n1478), .Y(n2149) );
  AO22X1_RVT U1460 ( .A1(n1151), .A2(n1516), .A3(n1147), .A4(n1152), .Y(N1051)
         );
  AO221X1_RVT U1461 ( .A1(N2536), .A2(n214), .A3(tmp_m1[22]), .A4(n213), .A5(
        N2801), .Y(n229) );
  INVX1_RVT U1462 ( .A(n1442), .Y(n1443) );
  INVX1_RVT U1463 ( .A(N1060), .Y(n1442) );
  OR3X2_RVT U1464 ( .A1(n2047), .A2(n2046), .A3(n2045), .Y(N1075) );
  INVX1_RVT U1465 ( .A(n1451), .Y(n1452) );
  INVX1_RVT U1466 ( .A(N1053), .Y(n1451) );
  INVX1_RVT U1467 ( .A(N1056), .Y(n1440) );
  NAND2X0_RVT U1468 ( .A1(n1444), .A2(n1445), .Y(N1057) );
  INVX1_RVT U1469 ( .A(n1735), .Y(N2055) );
  INVX1_RVT U1470 ( .A(n1433), .Y(n1431) );
  NAND2X0_RVT U1471 ( .A1(n1614), .A2(n1745), .Y(N2096) );
  NAND2X0_RVT U1472 ( .A1(n621), .A2(n622), .Y(n616) );
  AO221X1_RVT U1473 ( .A1(n583), .A2(n1850), .A3(tmp_m0[37]), .A4(n1857), .A5(
        n584), .Y(N2102) );
  NAND4X0_RVT U1474 ( .A1(n569), .A2(n570), .A3(n571), .A4(n1583), .Y(n567) );
  NOR2X1_RVT U1475 ( .A1(n535), .A2(n1689), .Y(n1714) );
  NOR2X1_RVT U1476 ( .A1(n510), .A2(n1693), .Y(n1729) );
  NAND3X0_RVT U1477 ( .A1(n1851), .A2(n1863), .A3(tmp_m0[0]), .Y(n2142) );
  INVX1_RVT U1478 ( .A(n1629), .Y(n1630) );
  INVX1_RVT U1479 ( .A(n1749), .Y(N2111) );
  AND2X1_RVT U1480 ( .A1(n1632), .A2(n1631), .Y(n1749) );
  AO221X1_RVT U1481 ( .A1(N248), .A2(net32930), .A3(N222), .A4(net27434), .A5(
        n2028), .Y(n2029) );
  NAND2X0_RVT U1482 ( .A1(n1453), .A2(n1454), .Y(N1054) );
  OR3X1_RVT U1483 ( .A1(n1412), .A2(n1413), .A3(n1414), .Y(N1055) );
  AO22X1_RVT U1484 ( .A1(N153), .A2(net32926), .A3(N462), .A4(net32958), .Y(
        n1412) );
  INVX1_RVT U1485 ( .A(net47575), .Y(net32926) );
  INVX1_RVT U1486 ( .A(net47614), .Y(net32958) );
  AO222X1_RVT U1487 ( .A1(N437), .A2(net32946), .A3(N353), .A4(net32952), .A5(
        N411), .A6(net32962), .Y(n1413) );
  INVX1_RVT U1488 ( .A(net32948), .Y(net32946) );
  INVX1_RVT U1489 ( .A(net47581), .Y(net32952) );
  INVX1_RVT U1490 ( .A(net27586), .Y(net32962) );
  AO221X1_RVT U1491 ( .A1(N237), .A2(net32932), .A3(N211), .A4(net32938), .A5(
        n1415), .Y(n1414) );
  INVX1_RVT U1492 ( .A(net36423), .Y(net32932) );
  INVX1_RVT U1493 ( .A(net27580), .Y(net32938) );
  AO22X1_RVT U1494 ( .A1(N997), .A2(net32880), .A3(N940), .A4(net32866), .Y(
        n1415) );
  INVX1_RVT U1495 ( .A(n1154), .Y(net32880) );
  INVX1_RVT U1496 ( .A(n1153), .Y(net32866) );
  NBUFFX2_RVT U1497 ( .A(n1657), .Y(n1417) );
  NBUFFX2_RVT U1498 ( .A(n1659), .Y(n1418) );
  INVX0_RVT U1499 ( .A(n1588), .Y(n1891) );
  NBUFFX2_RVT U1500 ( .A(n1649), .Y(n1419) );
  NBUFFX2_RVT U1501 ( .A(n1647), .Y(n1420) );
  NBUFFX2_RVT U1502 ( .A(n1653), .Y(n1421) );
  NBUFFX2_RVT U1503 ( .A(n1655), .Y(n1422) );
  NBUFFX2_RVT U1504 ( .A(n1651), .Y(n1423) );
  INVX1_RVT U1505 ( .A(n1424), .Y(n1425) );
  INVX0_RVT U1506 ( .A(n1697), .Y(n1817) );
  IBUFFX16_RVT U1507 ( .A(n1428), .Y(n1426) );
  IBUFFX16_RVT U1508 ( .A(n1426), .Y(n1427) );
  IBUFFX16_RVT U1509 ( .A(n1430), .Y(n1428) );
  IBUFFX4_RVT U1510 ( .A(n1438), .Y(n1702) );
  IBUFFX16_RVT U1511 ( .A(n1427), .Y(n1912) );
  INVX1_RVT U1512 ( .A(n1912), .Y(n1736) );
  AND2X1_RVT U1513 ( .A1(n1431), .A2(n1432), .Y(n1735) );
  NOR2X1_RVT U1514 ( .A1(n984), .A2(n1737), .Y(n1432) );
  NOR2X0_RVT U1515 ( .A1(n1534), .A2(n1434), .Y(n1584) );
  NAND2X0_RVT U1516 ( .A1(n1436), .A2(n987), .Y(n1434) );
  OR2X1_RVT U1517 ( .A1(n1750), .A2(n1751), .Y(n1435) );
  AND4X2_RVT U1518 ( .A1(n456), .A2(n457), .A3(n458), .A4(n459), .Y(n1626) );
  NOR3X0_RVT U1519 ( .A1(n1005), .A2(n1007), .A3(n1006), .Y(n1436) );
  OAI222X1_RVT U1520 ( .A1(n1912), .A2(n1818), .A3(n1912), .A4(n1805), .A5(
        n1736), .A6(n1702), .Y(n1534) );
  IBUFFX4_RVT U1521 ( .A(n1760), .Y(n1437) );
  INVX32_RVT U1522 ( .A(n1437), .Y(n1438) );
  NOR3X0_RVT U1523 ( .A1(n2112), .A2(n2111), .A3(n2110), .Y(N1056) );
  AOI221X1_RVT U1524 ( .A1(N962), .A2(net32866), .A3(N1019), .A4(net32876), 
        .A5(n1856), .Y(N1077) );
  INVX1_RVT U1525 ( .A(N1077), .Y(n1441) );
  OR3X2_RVT U1526 ( .A1(n2086), .A2(n2085), .A3(n2084), .Y(N1060) );
  INVX0_RVT U1527 ( .A(n2105), .Y(n1446) );
  INVX0_RVT U1528 ( .A(n2107), .Y(n1444) );
  NAND2X0_RVT U1529 ( .A1(n1446), .A2(n1447), .Y(n1448) );
  IBUFFX4_RVT U1530 ( .A(n1448), .Y(n1445) );
  INVX16_RVT U1531 ( .A(n1449), .Y(n1450) );
  OR3X1_RVT U1532 ( .A1(n2122), .A2(n2121), .A3(n2120), .Y(N1053) );
  INVX0_RVT U1533 ( .A(n2117), .Y(n1456) );
  INVX0_RVT U1534 ( .A(n2118), .Y(n1453) );
  NAND2X0_RVT U1535 ( .A1(n1455), .A2(n1456), .Y(n1457) );
  IBUFFX4_RVT U1536 ( .A(n1457), .Y(n1454) );
  AND3X1_RVT U1537 ( .A1(n330), .A2(n2487), .A3(N2450), .Y(n1463) );
  AND2X1_RVT U1538 ( .A1(tmp_m0[23]), .A2(n1844), .Y(n1471) );
  AND2X1_RVT U1539 ( .A1(tmp_m0[22]), .A2(n1699), .Y(n1477) );
  INVX0_RVT U1540 ( .A(n1867), .Y(n1871) );
  AOI222X1_RVT U1541 ( .A1(N1674), .A2(n1871), .A3(n1526), .A4(n1471), .A5(
        N1891), .A6(tmp_m0[24]), .Y(n1479) );
  INVX0_RVT U1542 ( .A(n1884), .Y(n1890) );
  AND3X1_RVT U1543 ( .A1(n1775), .A2(n1790), .A3(n2103), .Y(n1487) );
  AND3X1_RVT U1544 ( .A1(n1519), .A2(n1469), .A3(n1801), .Y(n1491) );
  INVX1_RVT U1545 ( .A(n580), .Y(n1820) );
  AOI222X1_RVT U1546 ( .A1(N1752), .A2(n1862), .A3(N1328), .A4(n1785), .A5(
        N1742), .A6(n1898), .Y(n1498) );
  AOI222X1_RVT U1547 ( .A1(N1751), .A2(n1862), .A3(N1327), .A4(n1785), .A5(
        N1741), .A6(n1897), .Y(n1499) );
  AOI222X1_RVT U1548 ( .A1(N1746), .A2(n1862), .A3(N1322), .A4(n1785), .A5(
        N1736), .A6(n1896), .Y(n1500) );
  AOI222X1_RVT U1549 ( .A1(N1747), .A2(n1862), .A3(N1323), .A4(n1785), .A5(
        N1737), .A6(n1896), .Y(n1501) );
  AOI222X1_RVT U1550 ( .A1(N1675), .A2(n1871), .A3(n1527), .A4(n1471), .A5(
        N1892), .A6(tmp_m0[24]), .Y(n1502) );
  AOI222X1_RVT U1551 ( .A1(N1676), .A2(n1871), .A3(n1525), .A4(n1471), .A5(
        N1893), .A6(tmp_m0[24]), .Y(n1503) );
  AND2X1_RVT U1552 ( .A1(n2102), .A2(n1473), .Y(n1519) );
  INVX1_RVT U1553 ( .A(tmp_m0[16]), .Y(n1842) );
  INVX1_RVT U1554 ( .A(n573), .Y(n1823) );
  AOI222X1_RVT U1555 ( .A1(N1748), .A2(n1862), .A3(N1324), .A4(n1785), .A5(
        N1738), .A6(n1896), .Y(n1521) );
  AOI222X1_RVT U1556 ( .A1(N1749), .A2(n1862), .A3(N1325), .A4(n1785), .A5(
        N1739), .A6(n1897), .Y(n1522) );
  AOI222X1_RVT U1557 ( .A1(N1750), .A2(n1862), .A3(N1326), .A4(n1785), .A5(
        N1740), .A6(n1897), .Y(n1523) );
  AOI222X1_RVT U1558 ( .A1(N1678), .A2(n1871), .A3(n1927), .A4(n1471), .A5(
        N1895), .A6(tmp_m0[24]), .Y(n1524) );
  AOI222X1_RVT U1559 ( .A1(N1662), .A2(n1882), .A3(N1812), .A4(n1888), .A5(
        N1822), .A6(n1477), .Y(n1529) );
  AOI222X1_RVT U1560 ( .A1(N1663), .A2(n1882), .A3(N1813), .A4(n1889), .A5(
        N1823), .A6(n1878), .Y(n1530) );
  AOI222X1_RVT U1561 ( .A1(N1667), .A2(n1882), .A3(N1817), .A4(n1889), .A5(
        N1827), .A6(n1878), .Y(n1531) );
  INVX0_RVT U1562 ( .A(n1765), .Y(n1825) );
  AO222X1_RVT U1563 ( .A1(tmp_m0[41]), .A2(n1863), .A3(n1785), .A4(tmp_m0[29]), 
        .A5(n1807), .A6(n503), .Y(n1532) );
  INVX1_RVT U1564 ( .A(n1491), .Y(n1802) );
  NAND2X0_RVT U1565 ( .A1(tmp_m0[20]), .A2(n1761), .Y(n1540) );
  OAI222X1_RVT U1566 ( .A1(n1797), .A2(net32948), .A3(n1798), .A4(net47581), 
        .A5(n1799), .A6(net27586), .Y(n1541) );
  AOI222X1_RVT U1567 ( .A1(N1661), .A2(n1882), .A3(N1811), .A4(n1888), .A5(
        N1821), .A6(n1477), .Y(n1542) );
  AND3X1_RVT U1568 ( .A1(tmp_m0[10]), .A2(n1519), .A3(n1801), .Y(n1543) );
  AND2X1_RVT U1569 ( .A1(tmp_m0[12]), .A2(n2102), .Y(n1544) );
  INVX1_RVT U1570 ( .A(n1487), .Y(n1822) );
  INVX1_RVT U1571 ( .A(n1774), .Y(n1819) );
  AOI222X1_RVT U1572 ( .A1(N1668), .A2(n1883), .A3(N1818), .A4(n1889), .A5(
        N1828), .A6(n1878), .Y(n1549) );
  AOI222X1_RVT U1573 ( .A1(N1664), .A2(n1882), .A3(N1814), .A4(n1889), .A5(
        N1824), .A6(n1878), .Y(n1550) );
  AOI222X1_RVT U1574 ( .A1(N1665), .A2(n1882), .A3(N1815), .A4(n1889), .A5(
        N1825), .A6(n1878), .Y(n1551) );
  AOI222X1_RVT U1575 ( .A1(N1666), .A2(n1882), .A3(N1816), .A4(n1889), .A5(
        N1826), .A6(n1878), .Y(n1552) );
  AOI222X1_RVT U1576 ( .A1(N1672), .A2(n1872), .A3(n1905), .A4(n1471), .A5(
        N1889), .A6(tmp_m0[24]), .Y(n1553) );
  AOI222X1_RVT U1577 ( .A1(N1673), .A2(n1872), .A3(n1916), .A4(n1471), .A5(
        N1890), .A6(tmp_m0[24]), .Y(n1554) );
  AOI222X1_RVT U1578 ( .A1(N1677), .A2(n1872), .A3(n1924), .A4(n1471), .A5(
        N1894), .A6(tmp_m0[24]), .Y(n1555) );
  INVX1_RVT U1579 ( .A(n1477), .Y(n1876) );
  OAI221X1_RVT U1580 ( .A1(n2316), .A2(n1805), .A3(n1475), .A4(n486), .A5(n502), .Y(n1556) );
  NAND2X0_RVT U1581 ( .A1(n328), .A2(n2483), .Y(n1557) );
  AND3X1_RVT U1582 ( .A1(n2458), .A2(n2474), .A3(n2441), .Y(n1558) );
  AOI221X1_RVT U1583 ( .A1(tmp_m0[28]), .A2(n1823), .A3(tmp_m0[27]), .A4(n2480), .A5(n1777), .Y(n1583) );
  INVX1_RVT U1584 ( .A(n2010), .Y(n1015) );
  NBUFFX2_RVT U1585 ( .A(n1793), .Y(n1824) );
  INVX1_RVT U1586 ( .A(n486), .Y(n1814) );
  AND2X1_RVT U1587 ( .A1(n1761), .A2(n1518), .Y(n1586) );
  AO221X1_RVT U1588 ( .A1(n2239), .A2(n1852), .A3(tmp_m0[17]), .A4(n1859), 
        .A5(n2238), .Y(n1587) );
  AND2X1_RVT U1589 ( .A1(tmp_m0[19]), .A2(n1586), .Y(n1588) );
  AO221X1_RVT U1590 ( .A1(n2248), .A2(n1851), .A3(tmp_m0[18]), .A4(n1859), 
        .A5(n2247), .Y(n1589) );
  AOI222X1_RVT U1591 ( .A1(tmp_m0[20]), .A2(tmp_m0[24]), .A3(n1765), .A4(
        tmp_m0[1]), .A5(n1425), .A6(tmp_m0[15]), .Y(n1590) );
  INVX1_RVT U1592 ( .A(n1544), .Y(n1821) );
  AND2X1_RVT U1593 ( .A1(n2315), .A2(n1497), .Y(n1593) );
  NAND2X0_RVT U1594 ( .A1(n2012), .A2(n1516), .Y(net47614) );
  AO221X1_RVT U1595 ( .A1(n2184), .A2(n1852), .A3(tmp_m0[11]), .A4(n1858), 
        .A5(n2183), .Y(n1596) );
  AOI222X1_RVT U1596 ( .A1(n1591), .A2(n1817), .A3(n1904), .A4(n2321), .A5(
        N1597), .A6(n1439), .Y(n1597) );
  AOI222X1_RVT U1597 ( .A1(N1588), .A2(n1817), .A3(n1592), .A4(n2321), .A5(
        N1598), .A6(n1439), .Y(n1598) );
  AOI222X1_RVT U1598 ( .A1(N1589), .A2(n1817), .A3(N1314), .A4(n2321), .A5(
        N1599), .A6(n1439), .Y(n1599) );
  AOI222X1_RVT U1599 ( .A1(N1590), .A2(n1817), .A3(N1315), .A4(n2321), .A5(
        N1600), .A6(n1439), .Y(n1600) );
  AOI222X1_RVT U1600 ( .A1(N1591), .A2(n1817), .A3(N1316), .A4(n2321), .A5(
        N1601), .A6(n1439), .Y(n1601) );
  AOI222X1_RVT U1601 ( .A1(N1592), .A2(n1817), .A3(N1317), .A4(n2321), .A5(
        N1602), .A6(n1439), .Y(n1602) );
  AOI222X1_RVT U1602 ( .A1(N1593), .A2(n1817), .A3(N1318), .A4(n2321), .A5(
        N1603), .A6(n1439), .Y(n1603) );
  INVX1_RVT U1603 ( .A(n1540), .Y(n1863) );
  INVX1_RVT U1604 ( .A(net27586), .Y(net27438) );
  AND4X1_RVT U1605 ( .A1(n418), .A2(n419), .A3(n420), .A4(n421), .Y(n1604) );
  INVX1_RVT U1606 ( .A(net27580), .Y(net27434) );
  AOI222X1_RVT U1607 ( .A1(N1671), .A2(n1872), .A3(n1908), .A4(n1471), .A5(
        N1888), .A6(tmp_m0[24]), .Y(n1607) );
  AOI22X1_RVT U1608 ( .A1(n1864), .A2(tmp_m0[32]), .A3(n1848), .A4(tmp_m0[30]), 
        .Y(n1614) );
  NAND3X0_RVT U1609 ( .A1(n454), .A2(sel_1[1]), .A3(n1585), .Y(n1616) );
  OR2X1_RVT U1610 ( .A1(sel_0[1]), .A2(n2014), .Y(net47581) );
  INVX1_RVT U1611 ( .A(n1853), .Y(n1850) );
  AOI22X1_RVT U1612 ( .A1(n1865), .A2(tmp_m0[35]), .A3(n1848), .A4(tmp_m0[33]), 
        .Y(n1618) );
  AOI22X1_RVT U1613 ( .A1(n1865), .A2(tmp_m0[37]), .A3(n1847), .A4(tmp_m0[35]), 
        .Y(n1619) );
  AO221X1_RVT U1614 ( .A1(n2192), .A2(n1852), .A3(tmp_m0[12]), .A4(n1858), 
        .A5(n2191), .Y(n1620) );
  AOI222X1_RVT U1615 ( .A1(n1908), .A2(n1817), .A3(n1908), .A4(n2321), .A5(
        N1596), .A6(n1439), .Y(n1621) );
  OR2X1_RVT U1616 ( .A1(sel_0[1]), .A2(n2011), .Y(net47575) );
  AO221X1_RVT U1617 ( .A1(n2180), .A2(n1852), .A3(tmp_m0[10]), .A4(n1858), 
        .A5(n2179), .Y(n1622) );
  OAI222X1_RVT U1618 ( .A1(n1476), .A2(n1868), .A3(n1625), .A4(n1844), .A5(
        n1795), .A6(n1873), .Y(n1624) );
  NAND4X1_RVT U1619 ( .A1(n2284), .A2(n2283), .A3(n2282), .A4(n2281), .Y(n2286) );
  NAND4X1_RVT U1620 ( .A1(n2218), .A2(n2217), .A3(n2216), .A4(n2215), .Y(n2220) );
  NAND4X1_RVT U1621 ( .A1(n2229), .A2(n2228), .A3(n2227), .A4(n2226), .Y(n2231) );
  NAND4X1_RVT U1622 ( .A1(n547), .A2(n548), .A3(n549), .A4(n550), .Y(n545) );
  IBUFFX4_RVT U1623 ( .A(n1620), .Y(n1627) );
  INVX1_RVT U1624 ( .A(n1627), .Y(n1628) );
  INVX1_RVT U1625 ( .A(N2111), .Y(n1629) );
  AOI21X1_RVT U1626 ( .A1(tmp_m0[46]), .A2(n452), .A3(n1865), .Y(n1632) );
  NAND4X0_RVT U1627 ( .A1(n1597), .A2(n1500), .A3(n1529), .A4(n1553), .Y(n1647) );
  OR4X1_RVT U1628 ( .A1(n948), .A2(n949), .A3(n950), .A4(n951), .Y(n1648) );
  NAND4X0_RVT U1629 ( .A1(n1598), .A2(n1501), .A3(n1530), .A4(n1554), .Y(n1649) );
  OR4X1_RVT U1630 ( .A1(n935), .A2(n936), .A3(n937), .A4(n938), .Y(n1650) );
  NAND4X0_RVT U1631 ( .A1(n1599), .A2(n1521), .A3(n1550), .A4(n1479), .Y(n1651) );
  OR4X1_RVT U1632 ( .A1(n922), .A2(n923), .A3(n924), .A4(n925), .Y(n1652) );
  NAND4X0_RVT U1633 ( .A1(n1600), .A2(n1522), .A3(n1551), .A4(n1502), .Y(n1653) );
  OR4X1_RVT U1634 ( .A1(n909), .A2(n910), .A3(n911), .A4(n912), .Y(n1654) );
  NAND4X0_RVT U1635 ( .A1(n1601), .A2(n1523), .A3(n1552), .A4(n1503), .Y(n1655) );
  OR4X1_RVT U1636 ( .A1(n896), .A2(n897), .A3(n898), .A4(n899), .Y(n1656) );
  NAND4X0_RVT U1637 ( .A1(n1602), .A2(n1499), .A3(n1531), .A4(n1555), .Y(n1657) );
  OR4X1_RVT U1638 ( .A1(n883), .A2(n884), .A3(n885), .A4(n886), .Y(n1658) );
  INVX1_RVT U1639 ( .A(n648), .Y(n1807) );
  INVX1_RVT U1640 ( .A(n1808), .Y(n2320) );
  NAND4X0_RVT U1641 ( .A1(n1603), .A2(n1498), .A3(n1549), .A4(n1524), .Y(n1659) );
  OR4X1_RVT U1642 ( .A1(n855), .A2(n856), .A3(n857), .A4(n858), .Y(n1660) );
  IBUFFX32_RVT U1643 ( .A(n2196), .Y(n1661) );
  IBUFFX32_RVT U1644 ( .A(n1721), .Y(N2107) );
  NOR2X1_RVT U1645 ( .A1(n1853), .A2(n1626), .Y(n1751) );
  AND2X1_RVT U1646 ( .A1(n2108), .A2(n2322), .Y(n1765) );
  OR4X1_RVT U1647 ( .A1(n1662), .A2(n1663), .A3(n1664), .A4(n1661), .Y(n2198)
         );
  OAI221X1_RVT U1648 ( .A1(n1860), .A2(n1469), .A3(n1702), .A4(n1494), .A5(
        n2193), .Y(n1662) );
  OAI221X1_RVT U1649 ( .A1(n1877), .A2(n1473), .A3(n1880), .A4(n1813), .A5(
        n2194), .Y(n1663) );
  OAI221X1_RVT U1650 ( .A1(n577), .A2(n2289), .A3(n576), .A4(n1533), .A5(n2195), .Y(n1664) );
  OR4X1_RVT U1651 ( .A1(n1666), .A2(n1667), .A3(n1668), .A4(n1665), .Y(n2271)
         );
  OAI221X1_RVT U1652 ( .A1(n1874), .A2(n1518), .A3(n1861), .A4(n1468), .A5(
        n2267), .Y(n1667) );
  OAI221X1_RVT U1653 ( .A1(n1887), .A2(n1484), .A3(n1875), .A4(n1492), .A5(
        n2268), .Y(n1668) );
  INVX8_RVT U1654 ( .A(n1929), .Y(n1928) );
  OR4X1_RVT U1655 ( .A1(n1670), .A2(n1671), .A3(n1672), .A4(n1669), .Y(n2239)
         );
  OAI222X1_RVT U1656 ( .A1(n1874), .A2(n1468), .A3(n1815), .A4(n1533), .A5(
        n1861), .A6(n1790), .Y(n1671) );
  OAI222X1_RVT U1657 ( .A1(n1876), .A2(n1842), .A3(n1868), .A4(n1473), .A5(
        n1879), .A6(n1801), .Y(n1672) );
  OR4X1_RVT U1658 ( .A1(n1674), .A2(n1675), .A3(n1676), .A4(n1673), .Y(n2184)
         );
  OAI221X1_RVT U1659 ( .A1(n1860), .A2(n2301), .A3(n1702), .A4(n1497), .A5(
        n2181), .Y(n1674) );
  OAI222X1_RVT U1660 ( .A1(n1886), .A2(n1803), .A3(n1880), .A4(n1485), .A5(
        n1875), .A6(n1469), .Y(n1675) );
  OAI222X1_RVT U1661 ( .A1(n573), .A2(n1462), .A3(n1818), .A4(n2291), .A5(n574), .A6(n1533), .Y(n1676) );
  OR4X1_RVT U1662 ( .A1(n1678), .A2(n1679), .A3(n1680), .A4(n1677), .Y(n2180)
         );
  OAI222X1_RVT U1663 ( .A1(n1874), .A2(n1469), .A3(n1702), .A4(n2291), .A5(
        n1861), .A6(n1813), .Y(n1678) );
  OAI222X1_RVT U1664 ( .A1(n1876), .A2(n1803), .A3(n1868), .A4(n1485), .A5(
        n1879), .A6(n1497), .Y(n1679) );
  OAI222X1_RVT U1665 ( .A1(n573), .A2(n1533), .A3(n1885), .A4(n2301), .A5(
        n1818), .A6(n2287), .Y(n1680) );
  OR4X1_RVT U1666 ( .A1(n1682), .A2(n1683), .A3(n1684), .A4(n1681), .Y(n2248)
         );
  OAI222X1_RVT U1667 ( .A1(n1869), .A2(n1613), .A3(n1861), .A4(n1791), .A5(
        n1873), .A6(n1484), .Y(n1683) );
  OAI222X1_RVT U1668 ( .A1(n1886), .A2(n1842), .A3(n1880), .A4(n1473), .A5(
        n1875), .A6(n1468), .Y(n1684) );
  IBUFFX32_RVT U1669 ( .A(n1738), .Y(N2109) );
  NAND4X0_RVT U1670 ( .A1(n2190), .A2(n2189), .A3(n2188), .A4(n2187), .Y(n2192) );
  INVX4_RVT U1671 ( .A(n1727), .Y(n1685) );
  IBUFFX4_RVT U1672 ( .A(n1705), .Y(n1687) );
  INVX1_RVT U1673 ( .A(n1687), .Y(n1688) );
  NBUFFX32_RVT U1674 ( .A(n1718), .Y(n1689) );
  IBUFFX16_RVT U1675 ( .A(n1726), .Y(n1725) );
  IBUFFX16_RVT U1676 ( .A(N2110), .Y(n1705) );
  INVX4_RVT U1677 ( .A(n1810), .Y(n2319) );
  NBUFFX32_RVT U1678 ( .A(n1733), .Y(n1693) );
  IBUFFX16_RVT U1679 ( .A(n1701), .Y(n1696) );
  IBUFFX16_RVT U1680 ( .A(n1696), .Y(n1697) );
  IBUFFX8_RVT U1681 ( .A(n1700), .Y(n1701) );
  NOR4X1_RVT U1682 ( .A1(n979), .A2(n980), .A3(n981), .A4(n982), .Y(n972) );
  NAND4X0_RVT U1683 ( .A1(n482), .A2(n483), .A3(n484), .A4(n485), .Y(n479) );
  IBUFFX16_RVT U1684 ( .A(n1743), .Y(n1742) );
  INVX16_RVT U1685 ( .A(n1703), .Y(n1704) );
  AOI221X2_RVT U1686 ( .A1(n479), .A2(n1849), .A3(tmp_m0[45]), .A4(n1858), 
        .A5(n481), .Y(N2110) );
  NAND2X0_RVT U1687 ( .A1(n1618), .A2(n1706), .Y(N2099) );
  NAND2X0_RVT U1688 ( .A1(tmp_m0[34]), .A2(n1857), .Y(n1707) );
  NAND2X0_RVT U1689 ( .A1(n604), .A2(n1850), .Y(n1708) );
  NAND2X0_RVT U1690 ( .A1(n1707), .A2(n1708), .Y(n1709) );
  IBUFFX4_RVT U1691 ( .A(n1709), .Y(n1706) );
  NAND2X0_RVT U1692 ( .A1(n1619), .A2(n1710), .Y(N2101) );
  NAND2X0_RVT U1693 ( .A1(tmp_m0[36]), .A2(n1857), .Y(n1711) );
  NAND2X0_RVT U1694 ( .A1(n591), .A2(n1850), .Y(n1712) );
  NAND2X0_RVT U1695 ( .A1(n1711), .A2(n1712), .Y(n1713) );
  IBUFFX4_RVT U1696 ( .A(n1713), .Y(n1710) );
  INVX0_RVT U1697 ( .A(n1714), .Y(N2106) );
  NOR2X0_RVT U1698 ( .A1(n1770), .A2(n1612), .Y(n1716) );
  NOR2X4_RVT U1699 ( .A1(n1853), .A2(n1715), .Y(n1717) );
  NOR2X0_RVT U1700 ( .A1(n1716), .A2(n1717), .Y(n1719) );
  IBUFFX32_RVT U1701 ( .A(n1719), .Y(n1718) );
  AOI221X1_RVT U1702 ( .A1(n629), .A2(n1851), .A3(tmp_m0[29]), .A4(n617), .A5(
        n630), .Y(N2095) );
  INVX1_RVT U1703 ( .A(N2095), .Y(n1720) );
  IBUFFX32_RVT U1704 ( .A(n523), .Y(n1722) );
  NOR2X0_RVT U1705 ( .A1(n1770), .A2(n1611), .Y(n1723) );
  NOR2X4_RVT U1706 ( .A1(n1853), .A2(n1722), .Y(n1724) );
  NOR2X0_RVT U1707 ( .A1(n524), .A2(n1725), .Y(n1721) );
  NOR2X0_RVT U1708 ( .A1(n1723), .A2(n1724), .Y(n1726) );
  AO22X1_RVT U1709 ( .A1(n1865), .A2(tmp_m0[43]), .A3(n1847), .A4(tmp_m0[41]), 
        .Y(n524) );
  IBUFFX4_RVT U1710 ( .A(N2056), .Y(n1727) );
  INVX0_RVT U1711 ( .A(n1729), .Y(N2108) );
  NOR2X0_RVT U1712 ( .A1(n1770), .A2(n1615), .Y(n1731) );
  NOR2X4_RVT U1713 ( .A1(n1853), .A2(n1730), .Y(n1732) );
  NOR2X0_RVT U1714 ( .A1(n1731), .A2(n1732), .Y(n1734) );
  IBUFFX32_RVT U1715 ( .A(n1734), .Y(n1733) );
  NOR2X0_RVT U1716 ( .A1(n455), .A2(N1129), .Y(n1737) );
  NOR2X0_RVT U1717 ( .A1(n1770), .A2(n1795), .Y(n1740) );
  NOR2X0_RVT U1718 ( .A1(n496), .A2(n1742), .Y(n1738) );
  NOR2X1_RVT U1719 ( .A1(n1740), .A2(n1741), .Y(n1743) );
  AO22X1_RVT U1720 ( .A1(n1865), .A2(tmp_m0[45]), .A3(n1847), .A4(tmp_m0[43]), 
        .Y(n496) );
  AOI221X1_RVT U1721 ( .A1(n2148), .A2(n1852), .A3(tmp_m0[6]), .A4(n619), .A5(
        n2147), .Y(N2070) );
  INVX1_RVT U1722 ( .A(N2070), .Y(n1744) );
  NAND2X0_RVT U1723 ( .A1(tmp_m0[31]), .A2(n1857), .Y(n1746) );
  NAND2X0_RVT U1724 ( .A1(n623), .A2(n1851), .Y(n1747) );
  NAND2X0_RVT U1725 ( .A1(n1746), .A2(n1747), .Y(n1748) );
  IBUFFX4_RVT U1726 ( .A(n1748), .Y(n1745) );
  NOR2X0_RVT U1727 ( .A1(n1625), .A2(n1616), .Y(n1750) );
  INVX4_RVT U1728 ( .A(n1805), .Y(n2321) );
  AND3X1_RVT U1729 ( .A1(n1607), .A2(n1542), .A3(n1759), .Y(n1754) );
  AND2X1_RVT U1730 ( .A1(n1621), .A2(n1754), .Y(n1758) );
  NAND2X0_RVT U1731 ( .A1(n1758), .A2(n1757), .Y(n958) );
  INVX0_RVT U1732 ( .A(n1770), .Y(n1859) );
  INVX1_RVT U1733 ( .A(n2090), .Y(n1761) );
  IBUFFX4_RVT U1734 ( .A(n1809), .Y(n1810) );
  INVX1_RVT U1735 ( .A(n1424), .Y(n1895) );
  NAND2X0_RVT U1736 ( .A1(n2088), .A2(n994), .Y(n648) );
  INVX1_RVT U1737 ( .A(tmp_m0[24]), .Y(n1843) );
  NBUFFX2_RVT U1738 ( .A(n2302), .Y(n1803) );
  OA22X1_RVT U1739 ( .A1(n1802), .A2(n1504), .A3(n1545), .A4(n408), .Y(n521)
         );
  OA22X1_RVT U1740 ( .A1(n1802), .A2(n2316), .A3(n1690), .A4(n408), .Y(n532)
         );
  OA22X1_RVT U1741 ( .A1(n1802), .A2(n1486), .A3(n1623), .A4(n408), .Y(n472)
         );
  OA22X1_RVT U1742 ( .A1(n1802), .A2(n1545), .A3(n1470), .A4(n408), .Y(n492)
         );
  OA22X1_RVT U1743 ( .A1(n1802), .A2(n1690), .A3(n1486), .A4(n408), .Y(n506)
         );
  AND2X1_RVT U1744 ( .A1(tmp_m0[16]), .A2(n2320), .Y(n1760) );
  INVX0_RVT U1745 ( .A(n1890), .Y(n1887) );
  INVX0_RVT U1746 ( .A(n1883), .Y(n1880) );
  INVX0_RVT U1747 ( .A(n1878), .Y(n1875) );
  INVX0_RVT U1748 ( .A(n1871), .Y(n1869) );
  INVX0_RVT U1749 ( .A(n1871), .Y(n1870) );
  OR3X1_RVT U1750 ( .A1(n1755), .A2(n1756), .A3(n2027), .Y(N1065) );
  AO22X1_RVT U1751 ( .A1(N163), .A2(net32924), .A3(N472), .A4(net32956), .Y(
        n1755) );
  AO222X1_RVT U1752 ( .A1(N447), .A2(net27435), .A3(N363), .A4(net32950), .A5(
        N421), .A6(net32962), .Y(n1756) );
  INVX0_RVT U1753 ( .A(n1770), .Y(n1858) );
  INVX1_RVT U1754 ( .A(n1154), .Y(net32882) );
  INVX1_RVT U1755 ( .A(n2103), .Y(n2102) );
  NOR4X1_RVT U1756 ( .A1(n961), .A2(n962), .A3(n963), .A4(n964), .Y(n1757) );
  INVX1_RVT U1757 ( .A(n1616), .Y(n1847) );
  INVX1_RVT U1758 ( .A(N414), .Y(n1799) );
  INVX1_RVT U1759 ( .A(N356), .Y(n1798) );
  INVX0_RVT U1760 ( .A(n1780), .Y(n1866) );
  INVX0_RVT U1761 ( .A(n1780), .Y(n1864) );
  AND2X1_RVT U1762 ( .A1(tmp_m0[14]), .A2(n1775), .Y(n1774) );
  INVX2_RVT U1763 ( .A(b_m[0]), .Y(n1929) );
  INVX1_RVT U1764 ( .A(n1416), .Y(n1931) );
  INVX1_RVT U1765 ( .A(n1939), .Y(n1938) );
  INVX1_RVT U1766 ( .A(b_m[21]), .Y(n1939) );
  INVX1_RVT U1767 ( .A(n1937), .Y(n1936) );
  INVX1_RVT U1768 ( .A(b_m[17]), .Y(n1937) );
  INVX1_RVT U1769 ( .A(n1935), .Y(n1934) );
  INVX1_RVT U1770 ( .A(b_m[16]), .Y(n1935) );
  INVX1_RVT U1771 ( .A(b_m[8]), .Y(n1933) );
  OA21X1_RVT U1772 ( .A1(n2016), .A2(n2324), .A3(n2326), .Y(n2017) );
  INVX1_RVT U1773 ( .A(net27435), .Y(net32948) );
  INVX1_RVT U1774 ( .A(n1888), .Y(n1886) );
  INVX1_RVT U1775 ( .A(n2139), .Y(n2153) );
  INVX1_RVT U1776 ( .A(n1495), .Y(n1883) );
  INVX1_RVT U1777 ( .A(n574), .Y(n2480) );
  INVX1_RVT U1778 ( .A(n1153), .Y(net32864) );
  INVX1_RVT U1779 ( .A(n1882), .Y(n1881) );
  INVX1_RVT U1780 ( .A(n1495), .Y(n1882) );
  INVX1_RVT U1781 ( .A(n2330), .Y(n2338) );
  INVX1_RVT U1782 ( .A(n2329), .Y(n2337) );
  INVX1_RVT U1783 ( .A(n2328), .Y(n2336) );
  INVX0_RVT U1784 ( .A(n2331), .Y(n2339) );
  INVX0_RVT U1785 ( .A(n2332), .Y(n2340) );
  AO21X1_RVT U1786 ( .A1(N984), .A2(net32870), .A3(n1856), .Y(N1099) );
  INVX1_RVT U1787 ( .A(n1884), .Y(n1888) );
  INVX1_RVT U1788 ( .A(n1884), .Y(n1889) );
  INVX1_RVT U1789 ( .A(n1153), .Y(net32870) );
  INVX1_RVT U1790 ( .A(n1153), .Y(net32868) );
  INVX1_RVT U1791 ( .A(n180), .Y(n1854) );
  INVX1_RVT U1792 ( .A(n180), .Y(n1855) );
  AND2X1_RVT U1793 ( .A1(n2320), .A2(n1491), .Y(n867) );
  IBUFFX4_RVT U1794 ( .A(n1804), .Y(n1805) );
  INVX1_RVT U1795 ( .A(n1814), .Y(n1815) );
  NAND3X0_RVT U1796 ( .A1(n1762), .A2(n1763), .A3(n1764), .Y(N1068) );
  AOI22X1_RVT U1797 ( .A1(N166), .A2(net32926), .A3(N475), .A4(net32956), .Y(
        n1762) );
  AOI222X1_RVT U1798 ( .A1(N450), .A2(net27435), .A3(N366), .A4(net32950), 
        .A5(N424), .A6(net32962), .Y(n1763) );
  AOI221X1_RVT U1799 ( .A1(N250), .A2(net32932), .A3(N224), .A4(net32938), 
        .A5(n2021), .Y(n1764) );
  INVX1_RVT U1800 ( .A(n576), .Y(n2478) );
  AO221X1_RVT U1801 ( .A1(N1382), .A2(n867), .A3(N1141), .A4(n1800), .A5(n965), 
        .Y(n961) );
  AO22X1_RVT U1802 ( .A1(N1117), .A2(n870), .A3(N1131), .A4(n871), .Y(n965) );
  AO221X1_RVT U1803 ( .A1(N1383), .A2(n867), .A3(N1142), .A4(n1800), .A5(n952), 
        .Y(n948) );
  AO22X1_RVT U1804 ( .A1(N1118), .A2(n870), .A3(N1132), .A4(n871), .Y(n952) );
  AO221X1_RVT U1805 ( .A1(N1384), .A2(n867), .A3(N1143), .A4(n1800), .A5(n939), 
        .Y(n935) );
  AO22X1_RVT U1806 ( .A1(N1119), .A2(n870), .A3(N1133), .A4(n871), .Y(n939) );
  AO221X1_RVT U1807 ( .A1(N1385), .A2(n867), .A3(N1144), .A4(n1800), .A5(n926), 
        .Y(n922) );
  AO22X1_RVT U1808 ( .A1(N1120), .A2(n870), .A3(N1134), .A4(n871), .Y(n926) );
  AO221X1_RVT U1809 ( .A1(N1386), .A2(n867), .A3(N1145), .A4(n1800), .A5(n913), 
        .Y(n909) );
  AO22X1_RVT U1810 ( .A1(N1121), .A2(n870), .A3(N1135), .A4(n871), .Y(n913) );
  AO221X1_RVT U1811 ( .A1(N1387), .A2(n867), .A3(N1146), .A4(n1800), .A5(n900), 
        .Y(n896) );
  AO22X1_RVT U1812 ( .A1(N1122), .A2(n870), .A3(N1136), .A4(n871), .Y(n900) );
  AO221X1_RVT U1813 ( .A1(N1388), .A2(n867), .A3(N1147), .A4(n1800), .A5(n887), 
        .Y(n883) );
  AO22X1_RVT U1814 ( .A1(N1123), .A2(n870), .A3(N1137), .A4(n871), .Y(n887) );
  AO221X1_RVT U1815 ( .A1(N1389), .A2(n867), .A3(N1148), .A4(n1800), .A5(n869), 
        .Y(n855) );
  AO22X1_RVT U1816 ( .A1(N1124), .A2(n870), .A3(N1138), .A4(n871), .Y(n869) );
  AND2X1_RVT U1817 ( .A1(n2124), .A2(n2322), .Y(n1800) );
  AO221X1_RVT U1818 ( .A1(N1958), .A2(n1864), .A3(N2037), .A4(n2317), .A5(n957), .Y(N2057) );
  AO222X1_RVT U1819 ( .A1(N2047), .A2(n1845), .A3(n958), .A4(n1849), .A5(N1968), .A6(n2472), .Y(n957) );
  AO221X1_RVT U1820 ( .A1(N1959), .A2(n1864), .A3(N2038), .A4(n2317), .A5(n944), .Y(N2058) );
  AO222X1_RVT U1821 ( .A1(N2048), .A2(n1845), .A3(n945), .A4(n1849), .A5(N1969), .A6(n2472), .Y(n944) );
  AO221X1_RVT U1822 ( .A1(N1960), .A2(n1864), .A3(N2039), .A4(n2317), .A5(n931), .Y(N2059) );
  AO222X1_RVT U1823 ( .A1(N2049), .A2(n1845), .A3(n932), .A4(n1849), .A5(N1970), .A6(n2472), .Y(n931) );
  AO221X1_RVT U1824 ( .A1(N1961), .A2(n1864), .A3(N2040), .A4(n2317), .A5(n918), .Y(N2060) );
  AO222X1_RVT U1825 ( .A1(N2050), .A2(n1845), .A3(n919), .A4(n1849), .A5(N1971), .A6(n2472), .Y(n918) );
  AO221X1_RVT U1826 ( .A1(N1962), .A2(n1864), .A3(N2041), .A4(n2317), .A5(n905), .Y(N2061) );
  AO222X1_RVT U1827 ( .A1(N2051), .A2(n1845), .A3(n906), .A4(n1849), .A5(N1972), .A6(n2472), .Y(n905) );
  AO221X1_RVT U1828 ( .A1(N1963), .A2(n1864), .A3(N2042), .A4(n2317), .A5(n892), .Y(N2062) );
  AO222X1_RVT U1829 ( .A1(N2052), .A2(n1845), .A3(n893), .A4(n1849), .A5(N1973), .A6(n2472), .Y(n892) );
  AO221X1_RVT U1830 ( .A1(N1964), .A2(n1864), .A3(N2043), .A4(n2317), .A5(n879), .Y(N2063) );
  AO222X1_RVT U1831 ( .A1(N2053), .A2(n1845), .A3(n880), .A4(n1849), .A5(N1974), .A6(n2472), .Y(n879) );
  AO221X1_RVT U1832 ( .A1(N1965), .A2(n1864), .A3(N2044), .A4(n2317), .A5(n850), .Y(N2064) );
  AO222X1_RVT U1833 ( .A1(N2054), .A2(n1845), .A3(n851), .A4(n1849), .A5(N1975), .A6(n2472), .Y(n850) );
  NAND2X0_RVT U1834 ( .A1(n2124), .A2(n2322), .Y(n463) );
  AO222X1_RVT U1835 ( .A1(n1910), .A2(n2481), .A3(N1391), .A4(n2478), .A5(
        n1910), .A6(n2479), .Y(n975) );
  AO222X1_RVT U1836 ( .A1(N1190), .A2(n2481), .A3(N1393), .A4(n2478), .A5(
        N1449), .A6(n2479), .Y(n949) );
  AO222X1_RVT U1837 ( .A1(N1191), .A2(n2481), .A3(N1394), .A4(n2478), .A5(
        N1450), .A6(n2479), .Y(n936) );
  AO222X1_RVT U1838 ( .A1(N1192), .A2(n2481), .A3(N1395), .A4(n2478), .A5(
        N1451), .A6(n2479), .Y(n923) );
  AO222X1_RVT U1839 ( .A1(N1193), .A2(n2481), .A3(N1396), .A4(n2478), .A5(
        N1452), .A6(n2479), .Y(n910) );
  AO222X1_RVT U1840 ( .A1(N1194), .A2(n2481), .A3(N1397), .A4(n2478), .A5(
        N1453), .A6(n2479), .Y(n897) );
  AO222X1_RVT U1841 ( .A1(N1195), .A2(n2481), .A3(N1398), .A4(n2478), .A5(
        N1454), .A6(n2479), .Y(n884) );
  AO222X1_RVT U1842 ( .A1(N1196), .A2(n2481), .A3(N1399), .A4(n2478), .A5(
        N1455), .A6(n2479), .Y(n856) );
  INVX1_RVT U1843 ( .A(n1471), .Y(n1873) );
  INVX1_RVT U1844 ( .A(n1876), .Y(n1878) );
  INVX1_RVT U1845 ( .A(n1471), .Y(n1874) );
  NAND2X0_RVT U1846 ( .A1(n1544), .A2(n2320), .Y(n574) );
  INVX1_RVT U1847 ( .A(n1898), .Y(n1894) );
  INVX1_RVT U1848 ( .A(n1899), .Y(n1893) );
  AO222X1_RVT U1849 ( .A1(N1458), .A2(n2480), .A3(N1199), .A4(n2482), .A5(
        N1249), .A6(n1765), .Y(n963) );
  AO222X1_RVT U1850 ( .A1(N1459), .A2(n2480), .A3(N1200), .A4(n2482), .A5(
        N1250), .A6(n1765), .Y(n950) );
  AO222X1_RVT U1851 ( .A1(N1460), .A2(n2480), .A3(N1201), .A4(n2482), .A5(
        N1251), .A6(n1765), .Y(n937) );
  AO222X1_RVT U1852 ( .A1(N1461), .A2(n2480), .A3(N1202), .A4(n2482), .A5(
        N1252), .A6(n1765), .Y(n924) );
  AO222X1_RVT U1853 ( .A1(N1462), .A2(n2480), .A3(N1203), .A4(n2482), .A5(
        N1253), .A6(n1765), .Y(n911) );
  AO222X1_RVT U1854 ( .A1(N1463), .A2(n2480), .A3(N1204), .A4(n2482), .A5(
        N1254), .A6(n1765), .Y(n898) );
  AO222X1_RVT U1855 ( .A1(N1464), .A2(n2480), .A3(N1205), .A4(n2482), .A5(
        N1255), .A6(n1765), .Y(n885) );
  AO222X1_RVT U1856 ( .A1(N1465), .A2(n2480), .A3(N1206), .A4(n2482), .A5(
        N1256), .A6(n1765), .Y(n857) );
  INVX1_RVT U1857 ( .A(sel_1[1]), .Y(n1851) );
  INVX1_RVT U1858 ( .A(n1853), .Y(n1849) );
  INVX1_RVT U1859 ( .A(n1770), .Y(n1857) );
  INVX1_RVT U1860 ( .A(n1148), .Y(n2016) );
  INVX0_RVT U1861 ( .A(n1804), .Y(n1806) );
  AO222X1_RVT U1862 ( .A1(N1265), .A2(n1814), .A3(N1522), .A4(n1823), .A5(
        N1532), .A6(n1820), .Y(n886) );
  AO222X1_RVT U1863 ( .A1(N1264), .A2(n1814), .A3(N1521), .A4(n1823), .A5(
        N1531), .A6(n1820), .Y(n899) );
  AO222X1_RVT U1864 ( .A1(N1263), .A2(n1814), .A3(N1520), .A4(n1823), .A5(
        N1530), .A6(n1820), .Y(n912) );
  AO222X1_RVT U1865 ( .A1(N1262), .A2(n1814), .A3(N1519), .A4(n1823), .A5(
        N1529), .A6(n1820), .Y(n925) );
  AO222X1_RVT U1866 ( .A1(N1261), .A2(n1814), .A3(N1518), .A4(n1823), .A5(
        N1528), .A6(n1820), .Y(n938) );
  AO222X1_RVT U1867 ( .A1(N1260), .A2(n1814), .A3(N1517), .A4(n1823), .A5(
        N1527), .A6(n1820), .Y(n951) );
  AO222X1_RVT U1868 ( .A1(N1259), .A2(n1814), .A3(N1516), .A4(n1823), .A5(
        N1526), .A6(n1820), .Y(n964) );
  AO222X1_RVT U1869 ( .A1(N1266), .A2(n1814), .A3(N1523), .A4(n1823), .A5(
        N1533), .A6(n1820), .Y(n858) );
  INVX1_RVT U1870 ( .A(n1138), .Y(n2440) );
  INVX0_RVT U1871 ( .A(n1140), .Y(n2323) );
  AO222X1_RVT U1872 ( .A1(n1910), .A2(n1817), .A3(n1910), .A4(n2321), .A5(
        N1595), .A6(n1439), .Y(n979) );
  INVX1_RVT U1873 ( .A(n1853), .Y(n1852) );
  INVX1_RVT U1874 ( .A(n1870), .Y(n1872) );
  INVX1_RVT U1875 ( .A(n2010), .Y(n1856) );
  INVX1_RVT U1876 ( .A(n577), .Y(n2479) );
  INVX1_RVT U1877 ( .A(n343), .Y(n2444) );
  INVX1_RVT U1878 ( .A(n241), .Y(n2450) );
  INVX1_RVT U1879 ( .A(n157), .Y(n2445) );
  INVX1_RVT U1880 ( .A(n1826), .Y(n1829) );
  INVX1_RVT U1881 ( .A(n1557), .Y(n1832) );
  INVX1_RVT U1882 ( .A(n1557), .Y(n1831) );
  INVX1_RVT U1883 ( .A(n1557), .Y(n1830) );
  INVX1_RVT U1884 ( .A(n1826), .Y(n1828) );
  INVX1_RVT U1885 ( .A(n1826), .Y(n1827) );
  INVX1_RVT U1886 ( .A(n849), .Y(n2472) );
  AO21X1_RVT U1887 ( .A1(n1471), .A2(n1560), .A3(n1859), .Y(n620) );
  XNOR2X1_RVT U1888 ( .A1(n1927), .A2(n1766), .Y(N2054) );
  NAND2X0_RVT U1889 ( .A1(n1924), .A2(\add_489/carry[8] ), .Y(n1766) );
  INVX1_RVT U1890 ( .A(n167), .Y(n2441) );
  INVX1_RVT U1891 ( .A(n1771), .Y(n1838) );
  INVX1_RVT U1892 ( .A(n1862), .Y(n1861) );
  INVX1_RVT U1893 ( .A(n243), .Y(n2447) );
  INVX0_RVT U1894 ( .A(n1154), .Y(net32878) );
  INVX0_RVT U1895 ( .A(n1154), .Y(net32876) );
  INVX1_RVT U1896 ( .A(n1772), .Y(n1837) );
  INVX1_RVT U1897 ( .A(n1773), .Y(n1836) );
  INVX1_RVT U1898 ( .A(n464), .Y(n2481) );
  INVX1_RVT U1899 ( .A(net47614), .Y(net32956) );
  INVX1_RVT U1900 ( .A(n1948), .Y(n1960) );
  INVX1_RVT U1901 ( .A(n1948), .Y(n1958) );
  INVX1_RVT U1902 ( .A(n1948), .Y(n1962) );
  INVX1_RVT U1903 ( .A(n1948), .Y(n1970) );
  INVX1_RVT U1904 ( .A(n1948), .Y(n1972) );
  INVX1_RVT U1905 ( .A(n1948), .Y(n1966) );
  INVX1_RVT U1906 ( .A(n1948), .Y(n1964) );
  INVX1_RVT U1907 ( .A(n1947), .Y(n1961) );
  INVX1_RVT U1908 ( .A(n1947), .Y(n1959) );
  INVX1_RVT U1909 ( .A(n1947), .Y(n1968) );
  INVX1_RVT U1910 ( .A(n1947), .Y(n1969) );
  INVX1_RVT U1911 ( .A(n1947), .Y(n1967) );
  INVX1_RVT U1912 ( .A(n1947), .Y(n1965) );
  INVX1_RVT U1913 ( .A(n1947), .Y(n1963) );
  INVX1_RVT U1914 ( .A(n1947), .Y(n1974) );
  INVX1_RVT U1915 ( .A(n1947), .Y(n1957) );
  INVX1_RVT U1916 ( .A(n1948), .Y(n1976) );
  INVX1_RVT U1917 ( .A(n1947), .Y(n1977) );
  INVX1_RVT U1918 ( .A(n1946), .Y(n1971) );
  INVX1_RVT U1919 ( .A(n1946), .Y(n1973) );
  INVX1_RVT U1920 ( .A(n1947), .Y(n1978) );
  INVX1_RVT U1921 ( .A(n1946), .Y(n1975) );
  OA22X1_RVT U1922 ( .A1(n1486), .A2(n1822), .A3(n1470), .A4(n1819), .Y(n531)
         );
  OA22X1_RVT U1923 ( .A1(n1470), .A2(n1822), .A3(n1623), .A4(n1819), .Y(n520)
         );
  OA22X1_RVT U1924 ( .A1(n402), .A2(n1789), .A3(n1545), .A4(n1824), .Y(n507)
         );
  OA22X1_RVT U1925 ( .A1(n1623), .A2(n1822), .A3(n1787), .A4(n1819), .Y(n505)
         );
  INVX1_RVT U1926 ( .A(tmp_m0[24]), .Y(n1844) );
  OA22X1_RVT U1927 ( .A1(n402), .A2(n1520), .A3(n1824), .A4(n1470), .Y(n473)
         );
  OA22X1_RVT U1928 ( .A1(n1822), .A2(n1789), .A3(n1496), .A4(n1819), .Y(n471)
         );
  OA22X1_RVT U1929 ( .A1(n402), .A2(n1496), .A3(n1486), .A4(n1824), .Y(n493)
         );
  OA22X1_RVT U1930 ( .A1(n1787), .A2(n1822), .A3(n1819), .A4(n1789), .Y(n491)
         );
  AND2X1_RVT U1931 ( .A1(n2301), .A2(n1813), .Y(n1768) );
  INVX1_RVT U1932 ( .A(n1573), .Y(n1930) );
  INVX1_RVT U1933 ( .A(N440), .Y(n1797) );
  AO222X1_RVT U1934 ( .A1(N1744), .A2(n1862), .A3(N1320), .A4(n1812), .A5(
        n1910), .A6(n1895), .Y(n980) );
  AO222X1_RVT U1935 ( .A1(n1608), .A2(n1845), .A3(n971), .A4(n1849), .A5(N1967), .A6(n2472), .Y(n970) );
  AO222X1_RVT U1936 ( .A1(n1912), .A2(n1814), .A3(N1129), .A4(n1823), .A5(
        n1912), .A6(n1820), .Y(n991) );
  AO222X1_RVT U1937 ( .A1(N1129), .A2(n2481), .A3(n1912), .A4(n2478), .A5(
        N1129), .A6(n2479), .Y(n989) );
  AO222X1_RVT U1938 ( .A1(n1429), .A2(n2472), .A3(N1129), .A4(n1845), .A5(
        N1129), .A6(n1864), .Y(n984) );
  NOR2X1_RVT U1939 ( .A1(n994), .A2(n432), .Y(n871) );
  INVX1_RVT U1940 ( .A(n1610), .Y(n1907) );
  INVX1_RVT U1941 ( .A(n1592), .Y(n1915) );
  INVX1_RVT U1942 ( .A(n1591), .Y(n1904) );
  INVX1_RVT U1943 ( .A(n1591), .Y(n1903) );
  INVX1_RVT U1944 ( .A(n1592), .Y(n1914) );
  INVX1_RVT U1945 ( .A(n1610), .Y(n1908) );
  INVX1_RVT U1946 ( .A(n1595), .Y(n1925) );
  INVX1_RVT U1947 ( .A(n1608), .Y(n1910) );
  INVX1_RVT U1948 ( .A(n1594), .Y(n1924) );
  INVX1_RVT U1949 ( .A(n1591), .Y(n1902) );
  INVX1_RVT U1950 ( .A(n1546), .Y(n1917) );
  INVX1_RVT U1951 ( .A(n1547), .Y(n1919) );
  INVX1_RVT U1952 ( .A(n1548), .Y(n1921) );
  INVX1_RVT U1953 ( .A(n1546), .Y(n1918) );
  INVX1_RVT U1954 ( .A(n1547), .Y(n1920) );
  INVX1_RVT U1955 ( .A(n1548), .Y(n1922) );
  INVX1_RVT U1956 ( .A(n1595), .Y(n1926) );
  OA221X1_RVT U1957 ( .A1(n2316), .A2(n1825), .A3(n1475), .A4(n461), .A5(n462), 
        .Y(n459) );
  AO222X1_RVT U1958 ( .A1(n1610), .A2(n2481), .A3(N1392), .A4(n2478), .A5(
        n1610), .A6(n2479), .Y(n962) );
  OA221X1_RVT U1959 ( .A1(n1694), .A2(n1786), .A3(n1475), .A4(n1805), .A5(n516), .Y(n514) );
  AND3X1_RVT U1960 ( .A1(n1699), .A2(n1474), .A3(n2090), .Y(n1769) );
  OA221X1_RVT U1961 ( .A1(n2316), .A2(n1815), .A3(n1475), .A4(n1825), .A5(n487), .Y(n485) );
  OA221X1_RVT U1962 ( .A1(n1892), .A2(n1611), .A3(n1861), .A4(n1615), .A5(n475), .Y(n457) );
  OA22X1_RVT U1963 ( .A1(n1795), .A2(n1886), .A3(n1461), .A4(n1880), .Y(n475)
         );
  OA221X1_RVT U1964 ( .A1(n2316), .A2(n580), .A3(n1475), .A4(n573), .A5(n589), 
        .Y(n588) );
  OA22X1_RVT U1965 ( .A1(n1894), .A2(n1612), .A3(n1615), .A4(n1886), .Y(n494)
         );
  OA22X1_RVT U1966 ( .A1(n1461), .A2(n1893), .A3(n1885), .A4(n1611), .Y(n508)
         );
  OA221X1_RVT U1967 ( .A1(n2316), .A2(n1818), .A3(n1475), .A4(n580), .A5(n597), 
        .Y(n596) );
  AO222X1_RVT U1968 ( .A1(N1457), .A2(n2480), .A3(N1198), .A4(n2482), .A5(
        n1608), .A6(n1765), .Y(n976) );
  INVX1_RVT U1969 ( .A(n454), .Y(n2473) );
  INVX1_RVT U1970 ( .A(n1780), .Y(n1865) );
  AND2X1_RVT U1971 ( .A1(n849), .A2(n455), .Y(n1770) );
  OA22X1_RVT U1972 ( .A1(n1802), .A2(n1475), .A3(n1504), .A4(n408), .Y(n543)
         );
  OA22X1_RVT U1973 ( .A1(n402), .A2(n1470), .A3(n2316), .A4(n1824), .Y(n544)
         );
  INVX0_RVT U1974 ( .A(n2318), .Y(n1853) );
  OA22X1_RVT U1975 ( .A1(n1690), .A2(n1822), .A3(n1545), .A4(n1819), .Y(n553)
         );
  OA22X1_RVT U1976 ( .A1(n1545), .A2(n1822), .A3(n1486), .A4(n1819), .Y(n542)
         );
  OA22X1_RVT U1977 ( .A1(n402), .A2(n1476), .A3(n1824), .A4(n1623), .Y(n401)
         );
  OA22X1_RVT U1978 ( .A1(n1822), .A2(n1496), .A3(n1819), .A4(n1520), .Y(n399)
         );
  OA22X1_RVT U1979 ( .A1(n1802), .A2(n1470), .A3(n408), .A4(n1787), .Y(n400)
         );
  INVX1_RVT U1980 ( .A(n1616), .Y(n1845) );
  AND4X1_RVT U1981 ( .A1(n1761), .A2(n2315), .A3(n426), .A4(n428), .Y(n644) );
  INVX0_RVT U1982 ( .A(N94), .Y(n2439) );
  INVX1_RVT U1983 ( .A(N95), .Y(n2436) );
  INVX1_RVT U1984 ( .A(n1610), .Y(n1906) );
  INVX1_RVT U1985 ( .A(n1594), .Y(n1923) );
  INVX1_RVT U1986 ( .A(n1592), .Y(n1913) );
  AND2X1_RVT U1987 ( .A1(n2438), .A2(n1147), .Y(n1031) );
  INVX1_RVT U1988 ( .A(net47581), .Y(net32950) );
  OA22X1_RVT U1989 ( .A1(n1873), .A2(n1561), .A3(n1868), .A4(n1611), .Y(n389)
         );
  OR3X2_RVT U1990 ( .A1(n2004), .A2(N95), .A3(N94), .Y(n1148) );
  OA222X1_RVT U1991 ( .A1(n1461), .A2(n1874), .A3(n1623), .A4(n1881), .A5(
        n1476), .A6(n1875), .Y(n548) );
  OA222X1_RVT U1992 ( .A1(n1612), .A2(n1874), .A3(n1787), .A4(n1881), .A5(
        n1461), .A6(n1875), .Y(n537) );
  INVX1_RVT U1993 ( .A(net36423), .Y(net32930) );
  AO222X1_RVT U1994 ( .A1(N1258), .A2(n1814), .A3(n1608), .A4(n1823), .A5(
        N1525), .A6(n1820), .Y(n977) );
  INVX1_RVT U1995 ( .A(net47575), .Y(net32924) );
  OA22X1_RVT U1996 ( .A1(n1496), .A2(n1886), .A3(n1470), .A4(n1880), .Y(n560)
         );
  AND2X1_RVT U1997 ( .A1(n1162), .A2(n1516), .Y(n1165) );
  AO221X1_RVT U1998 ( .A1(N177), .A2(net32876), .A3(N929), .A4(net32868), .A5(
        n1171), .Y(N1042) );
  AO22X1_RVT U1999 ( .A1(n1164), .A2(b_e[1]), .A3(n1165), .A4(a_e[1]), .Y(
        n1171) );
  AO221X1_RVT U2000 ( .A1(N178), .A2(net32876), .A3(N930), .A4(net32868), .A5(
        n1170), .Y(N1043) );
  AO22X1_RVT U2001 ( .A1(n1164), .A2(b_e[2]), .A3(n1165), .A4(a_e[2]), .Y(
        n1170) );
  AO221X1_RVT U2002 ( .A1(N179), .A2(net32876), .A3(N931), .A4(net32864), .A5(
        n1169), .Y(N1044) );
  AO22X1_RVT U2003 ( .A1(n1164), .A2(b_e[3]), .A3(n1165), .A4(a_e[3]), .Y(
        n1169) );
  AO221X1_RVT U2004 ( .A1(N180), .A2(net32876), .A3(N932), .A4(net32868), .A5(
        n1168), .Y(N1045) );
  AO22X1_RVT U2005 ( .A1(n1164), .A2(b_e[4]), .A3(n1165), .A4(a_e[4]), .Y(
        n1168) );
  AO221X1_RVT U2006 ( .A1(N181), .A2(net32876), .A3(N933), .A4(net32870), .A5(
        n1167), .Y(N1046) );
  AO22X1_RVT U2007 ( .A1(n1164), .A2(b_e[5]), .A3(n1165), .A4(a_e[5]), .Y(
        n1167) );
  AO221X1_RVT U2008 ( .A1(N182), .A2(net32876), .A3(N934), .A4(net32870), .A5(
        n1166), .Y(N1047) );
  AO22X1_RVT U2009 ( .A1(n1164), .A2(b_e[6]), .A3(n1165), .A4(a_e[6]), .Y(
        n1166) );
  AO221X1_RVT U2010 ( .A1(N183), .A2(net32876), .A3(N935), .A4(net32870), .A5(
        n1163), .Y(N1048) );
  AO22X1_RVT U2011 ( .A1(n1164), .A2(b_e[7]), .A3(n1165), .A4(a_e[7]), .Y(
        n1163) );
  INVX1_RVT U2012 ( .A(n1616), .Y(n1846) );
  AO222X1_RVT U2013 ( .A1(n1608), .A2(n1882), .A3(n1608), .A4(n1888), .A5(
        N1820), .A6(n1477), .Y(n981) );
  INVX1_RVT U2014 ( .A(n2327), .Y(n2335) );
  OA222X1_RVT U2015 ( .A1(n1787), .A2(n1876), .A3(n1623), .A4(n1887), .A5(
        n1690), .A6(n1879), .Y(n594) );
  OA221X1_RVT U2016 ( .A1(n1789), .A2(n1876), .A3(n1545), .A4(n1880), .A5(n590), .Y(n586) );
  OA22X1_RVT U2017 ( .A1(n1470), .A2(n1893), .A3(n1787), .A4(n1886), .Y(n590)
         );
  AO222X1_RVT U2018 ( .A1(N1129), .A2(n1882), .A3(N1129), .A4(n1890), .A5(
        n1430), .A6(n1878), .Y(n1006) );
  INVX1_RVT U2019 ( .A(n1595), .Y(n1927) );
  INVX1_RVT U2020 ( .A(n1592), .Y(n1916) );
  INVX1_RVT U2021 ( .A(n1591), .Y(n1905) );
  OA221X1_RVT U2022 ( .A1(n1496), .A2(n1876), .A3(n1486), .A4(n1880), .A5(n582), .Y(n570) );
  OA22X1_RVT U2023 ( .A1(n1623), .A2(n1893), .A3(n1789), .A4(n1885), .Y(n582)
         );
  INVX1_RVT U2024 ( .A(n455), .Y(n2317) );
  OA222X1_RVT U2025 ( .A1(n1470), .A2(n1874), .A3(n1475), .A4(n1881), .A5(
        n1486), .A6(n1875), .Y(n613) );
  AO222X1_RVT U2026 ( .A1(n1912), .A2(n1862), .A3(n1430), .A4(n1809), .A5(
        N1129), .A6(n1895), .Y(n1005) );
  OA222X1_RVT U2027 ( .A1(n1623), .A2(n1874), .A3(n2316), .A4(n1881), .A5(
        n1470), .A6(n1875), .Y(n607) );
  OA222X1_RVT U2028 ( .A1(n1623), .A2(n1876), .A3(n1470), .A4(n1887), .A5(
        n1504), .A6(n1879), .Y(n601) );
  AND2X1_RVT U2029 ( .A1(n242), .A2(n172), .Y(n347) );
  INVX1_RVT U2030 ( .A(n156), .Y(n2448) );
  INVX1_RVT U2031 ( .A(n175), .Y(n2449) );
  INVX1_RVT U2032 ( .A(n169), .Y(n2465) );
  INVX1_RVT U2033 ( .A(n239), .Y(n2475) );
  INVX1_RVT U2034 ( .A(n214), .Y(n1826) );
  AND2X1_RVT U2035 ( .A1(n330), .A2(n2484), .Y(n214) );
  INVX1_RVT U2036 ( .A(N2450), .Y(n2484) );
  AO221X1_RVT U2037 ( .A1(n2475), .A2(n237), .A3(n2447), .A4(n2474), .A5(n223), 
        .Y(N2801) );
  OA22X1_RVT U2038 ( .A1(n167), .A2(n168), .A3(n169), .A4(n2447), .Y(n161) );
  AO221X1_RVT U2039 ( .A1(n339), .A2(n2474), .A3(n1854), .A4(n2458), .A5(n340), 
        .Y(N2768) );
  AO21X1_RVT U2040 ( .A1(N2233), .A2(n184), .A3(n2442), .Y(n340) );
  AO21X1_RVT U2041 ( .A1(n243), .A2(n167), .A3(n166), .Y(n339) );
  INVX1_RVT U2042 ( .A(n158), .Y(n2442) );
  INVX1_RVT U2043 ( .A(N2119), .Y(n2486) );
  AO22X1_RVT U2044 ( .A1(N2450), .A2(n330), .A3(N2230), .A4(n328), .Y(n184) );
  OA222X1_RVT U2045 ( .A1(n1486), .A2(n1886), .A3(n1545), .A4(n1860), .A5(
        n1690), .A6(n1892), .Y(n608) );
  OA22X1_RVT U2046 ( .A1(n1504), .A2(n1893), .A3(n1545), .A4(n1885), .Y(n614)
         );
  OA22X1_RVT U2047 ( .A1(n1690), .A2(n1876), .A3(n1545), .A4(n1874), .Y(n626)
         );
  OA22X1_RVT U2048 ( .A1(n1504), .A2(n580), .A3(n1690), .A4(n1818), .Y(n579)
         );
  INVX1_RVT U2049 ( .A(N2230), .Y(n2483) );
  INVX1_RVT U2050 ( .A(N2118), .Y(n2485) );
  INVX1_RVT U2051 ( .A(n1616), .Y(n1848) );
  OA222X1_RVT U2052 ( .A1(n1545), .A2(n1893), .A3(n2316), .A4(n1702), .A5(
        n1486), .A6(n1861), .Y(n602) );
  INVX1_RVT U2053 ( .A(n242), .Y(n2443) );
  AND2X1_RVT U2054 ( .A1(N993), .A2(net32876), .Y(N1050) );
  INVX1_RVT U2055 ( .A(n172), .Y(n2458) );
  AO21X1_RVT U2056 ( .A1(N936), .A2(net32870), .A3(N1050), .Y(N1049) );
  OA221X1_RVT U2057 ( .A1(n342), .A2(n239), .A3(n2474), .A4(n343), .A5(n344), 
        .Y(n158) );
  OA222X1_RVT U2058 ( .A1(n2443), .A2(n225), .A3(n347), .A4(n241), .A5(n2458), 
        .A6(n224), .Y(n342) );
  AO21X1_RVT U2059 ( .A1(n2443), .A2(n239), .A3(n346), .Y(n345) );
  INVX1_RVT U2060 ( .A(N2233), .Y(n2487) );
  INVX1_RVT U2061 ( .A(n1782), .Y(n1841) );
  INVX1_RVT U2062 ( .A(n1782), .Y(n1839) );
  INVX1_RVT U2063 ( .A(n1782), .Y(n1840) );
  OR2X1_RVT U2064 ( .A1(n2139), .A2(n2289), .Y(n2143) );
  OR2X1_RVT U2065 ( .A1(n2139), .A2(n1816), .Y(n2098) );
  OA22X1_RVT U2066 ( .A1(n173), .A2(n2447), .A3(n172), .A4(n167), .Y(n159) );
  OA21X1_RVT U2067 ( .A1(n2465), .A2(n164), .A3(n175), .Y(n173) );
  OA21X1_RVT U2068 ( .A1(n175), .A2(n169), .A3(n226), .Y(n243) );
  NAND3X0_RVT U2069 ( .A1(n330), .A2(n2487), .A3(N2450), .Y(n1771) );
  NAND3X0_RVT U2070 ( .A1(n328), .A2(n2487), .A3(N2230), .Y(n1772) );
  NAND3X0_RVT U2071 ( .A1(n328), .A2(n2487), .A3(N2230), .Y(n1773) );
  INVX1_RVT U2072 ( .A(n1558), .Y(n1833) );
  INVX0_RVT U2073 ( .A(n1143), .Y(n2005) );
  INVX1_RVT U2074 ( .A(n402), .Y(n2101) );
  INVX1_RVT U2075 ( .A(n1956), .Y(n1948) );
  INVX1_RVT U2076 ( .A(n1956), .Y(n1950) );
  INVX1_RVT U2077 ( .A(n1956), .Y(n1951) );
  INVX1_RVT U2078 ( .A(n1956), .Y(n1952) );
  INVX1_RVT U2079 ( .A(n1955), .Y(n1953) );
  INVX1_RVT U2080 ( .A(n1955), .Y(n1954) );
  INVX1_RVT U2081 ( .A(n1955), .Y(n1949) );
  INVX1_RVT U2082 ( .A(n1956), .Y(n1947) );
  INVX1_RVT U2083 ( .A(n1955), .Y(n1946) );
  INVX1_RVT U2084 ( .A(n1955), .Y(n1945) );
  INVX1_RVT U2085 ( .A(n1956), .Y(n1944) );
  INVX1_RVT U2086 ( .A(n1956), .Y(n1943) );
  INVX1_RVT U2087 ( .A(n1956), .Y(n1940) );
  INVX1_RVT U2088 ( .A(n1978), .Y(n1942) );
  INVX1_RVT U2089 ( .A(n1955), .Y(n1941) );
  OA222X1_RVT U2090 ( .A1(n1612), .A2(n1876), .A3(n1461), .A4(n1887), .A5(
        n1789), .A6(n1879), .Y(n526) );
  AO22X1_RVT U2091 ( .A1(n1865), .A2(tmp_m0[44]), .A3(n1847), .A4(tmp_m0[42]), 
        .Y(n510) );
  OA222X1_RVT U2092 ( .A1(n1877), .A2(n1611), .A3(n1885), .A4(n1612), .A5(
        n1496), .A6(n1879), .Y(n512) );
  OA22X1_RVT U2093 ( .A1(n402), .A2(n1623), .A3(n1504), .A4(n1824), .Y(n533)
         );
  OA22X1_RVT U2094 ( .A1(n402), .A2(n1787), .A3(n1690), .A4(n1824), .Y(n522)
         );
  AND2X1_RVT U2095 ( .A1(n1792), .A2(n1791), .Y(n1775) );
  OR4X1_RVT U2096 ( .A1(n1624), .A2(n1776), .A3(n1532), .A4(n1556), .Y(n495)
         );
  OAI221X1_RVT U2097 ( .A1(n1615), .A2(n1876), .A3(n1520), .A4(n1880), .A5(
        n508), .Y(n1776) );
  AOI221X1_RVT U2098 ( .A1(n1812), .A2(tmp_m0[31]), .A3(n1807), .A4(n466), 
        .A5(n467), .Y(n458) );
  AO22X1_RVT U2099 ( .A1(n2321), .A2(tmp_m0[30]), .A3(n1814), .A4(tmp_m0[29]), 
        .Y(n467) );
  AO22X1_RVT U2100 ( .A1(n2319), .A2(tmp_m0[30]), .A3(n2321), .A4(tmp_m0[29]), 
        .Y(n489) );
  AO22X1_RVT U2101 ( .A1(n1864), .A2(tmp_m0[46]), .A3(n1847), .A4(tmp_m0[44]), 
        .Y(n481) );
  OA221X1_RVT U2102 ( .A1(n1795), .A2(n1876), .A3(n1476), .A4(n1880), .A5(n494), .Y(n483) );
  AO22X1_RVT U2103 ( .A1(n2478), .A2(tmp_m0[25]), .A3(n2479), .A4(tmp_m0[26]), 
        .Y(n1777) );
  AO221X1_RVT U2104 ( .A1(n567), .A2(n1850), .A3(tmp_m0[38]), .A4(n1857), .A5(
        n568), .Y(N2103) );
  AO22X1_RVT U2105 ( .A1(n1865), .A2(tmp_m0[39]), .A3(n1847), .A4(tmp_m0[37]), 
        .Y(n568) );
  OA221X1_RVT U2106 ( .A1(n1787), .A2(n1860), .A3(n1545), .A4(n1702), .A5(n579), .Y(n571) );
  AO221X1_RVT U2107 ( .A1(n1608), .A2(n867), .A3(N1140), .A4(n1800), .A5(n978), 
        .Y(n974) );
  AO22X1_RVT U2108 ( .A1(N1116), .A2(n870), .A3(n1608), .A4(n871), .Y(n978) );
  OR2X1_RVT U2109 ( .A1(n2149), .A2(n1778), .Y(n2290) );
  AO221X1_RVT U2110 ( .A1(N1129), .A2(n867), .A3(n1912), .A4(n1800), .A5(n1000), .Y(n988) );
  AO22X1_RVT U2111 ( .A1(n1430), .A2(n870), .A3(N1129), .A4(n871), .Y(n1000)
         );
  AND2X1_RVT U2112 ( .A1(tmp_m0[18]), .A2(n2099), .Y(n1779) );
  AO22X1_RVT U2113 ( .A1(n1865), .A2(tmp_m0[38]), .A3(n1847), .A4(tmp_m0[36]), 
        .Y(n584) );
  OA222X1_RVT U2114 ( .A1(n1623), .A2(n1860), .A3(n1504), .A4(n1818), .A5(
        n1690), .A6(n1702), .Y(n587) );
  OA222X1_RVT U2115 ( .A1(n1486), .A2(n1892), .A3(n1504), .A4(n1702), .A5(
        n1470), .A6(n1861), .Y(n595) );
  OR2X1_RVT U2116 ( .A1(n1851), .A2(sel_1[0]), .Y(n454) );
  NAND2X0_RVT U2117 ( .A1(n2473), .A2(tmp_m0[47]), .Y(n1780) );
  AO22X1_RVT U2118 ( .A1(n1865), .A2(tmp_m0[42]), .A3(n1847), .A4(tmp_m0[40]), 
        .Y(n535) );
  OA222X1_RVT U2119 ( .A1(n1476), .A2(n1886), .A3(n1520), .A4(n1860), .A5(
        n1496), .A6(n1892), .Y(n538) );
  AO222X1_RVT U2120 ( .A1(n1845), .A2(tmp_m0[46]), .A3(n386), .A4(n1849), .A5(
        n2317), .A6(tmp_m0[47]), .Y(N2112) );
  OA22X1_RVT U2121 ( .A1(n1894), .A2(n1615), .A3(n1885), .A4(n1625), .Y(n391)
         );
  OA22X1_RVT U2122 ( .A1(n1881), .A2(n1612), .A3(n1875), .A4(n1606), .Y(n390)
         );
  OA22X1_RVT U2123 ( .A1(n1486), .A2(n402), .A3(n1475), .A4(n1824), .Y(n555)
         );
  AO221X1_RVT U2124 ( .A1(n545), .A2(n1850), .A3(tmp_m0[40]), .A4(n1857), .A5(
        n546), .Y(N2105) );
  AO22X1_RVT U2125 ( .A1(n1865), .A2(tmp_m0[41]), .A3(n1847), .A4(tmp_m0[39]), 
        .Y(n546) );
  OA22X1_RVT U2126 ( .A1(n1789), .A2(n1893), .A3(n1520), .A4(n1886), .Y(n549)
         );
  AO22X1_RVT U2127 ( .A1(n1865), .A2(tmp_m0[40]), .A3(n1847), .A4(tmp_m0[38]), 
        .Y(n557) );
  OA22X1_RVT U2128 ( .A1(n1520), .A2(n1876), .A3(n1476), .A4(n1873), .Y(n559)
         );
  AND2X1_RVT U2129 ( .A1(sel_0[0]), .A2(n2326), .Y(n1781) );
  OA21X1_RVT U2130 ( .A1(n1138), .A2(sel_0[0]), .A3(n1139), .Y(n2014) );
  INVX0_RVT U2131 ( .A(n2368), .Y(n2370) );
  INVX0_RVT U2132 ( .A(n1162), .Y(n2437) );
  AO221X1_RVT U2133 ( .A1(n1398), .A2(n1155), .A3(n1156), .A4(n1605), .A5(
        n1157), .Y(n1151) );
  NAND2X0_RVT U2134 ( .A1(n2018), .A2(n1516), .Y(net36423) );
  OA21X1_RVT U2135 ( .A1(n1136), .A2(sel_0[0]), .A3(n1137), .Y(n2011) );
  OA22X1_RVT U2136 ( .A1(n2316), .A2(n1860), .A3(n1475), .A4(n1892), .Y(n628)
         );
  AO221X1_RVT U2137 ( .A1(n616), .A2(n1850), .A3(tmp_m0[31]), .A4(n617), .A5(
        n618), .Y(N2097) );
  AO22X1_RVT U2138 ( .A1(tmp_m0[33]), .A2(n619), .A3(tmp_m0[32]), .A4(n620), 
        .Y(n618) );
  AO22X1_RVT U2139 ( .A1(tmp_m0[31]), .A2(n619), .A3(tmp_m0[30]), .A4(n620), 
        .Y(n630) );
  AO221X1_RVT U2140 ( .A1(n598), .A2(n1850), .A3(tmp_m0[35]), .A4(n1857), .A5(
        n599), .Y(N2100) );
  AO22X1_RVT U2141 ( .A1(n1865), .A2(tmp_m0[36]), .A3(n1848), .A4(tmp_m0[34]), 
        .Y(n599) );
  AO221X1_RVT U2142 ( .A1(n610), .A2(n1851), .A3(tmp_m0[33]), .A4(n1857), .A5(
        n611), .Y(N2098) );
  AO22X1_RVT U2143 ( .A1(n1865), .A2(tmp_m0[34]), .A3(n1848), .A4(tmp_m0[32]), 
        .Y(n611) );
  AO221X1_RVT U2144 ( .A1(N176), .A2(net32876), .A3(N928), .A4(net32868), .A5(
        n1172), .Y(N1041) );
  AO22X1_RVT U2145 ( .A1(n1164), .A2(b_e[0]), .A3(n1165), .A4(a_e[0]), .Y(
        n1172) );
  AND2X1_RVT U2146 ( .A1(n1174), .A2(n1516), .Y(n1164) );
  AOI221X1_RVT U2147 ( .A1(n2474), .A2(n218), .A3(n2475), .A4(n220), .A5(n221), 
        .Y(n176) );
  AO221X1_RVT U2148 ( .A1(n2444), .A2(\sel_2[1] ), .A3(N2233), .A4(n184), .A5(
        n223), .Y(n221) );
  OA222X1_RVT U2149 ( .A1(n2384), .A2(n180), .A3(n181), .A4(n1178), .A5(n2457), 
        .A6(n1833), .Y(n210) );
  OA222X1_RVT U2150 ( .A1(n2385), .A2(n180), .A3(n181), .A4(n1179), .A5(n2456), 
        .A6(n1833), .Y(n206) );
  OA222X1_RVT U2151 ( .A1(n2470), .A2(n180), .A3(n181), .A4(n1180), .A5(n2455), 
        .A6(n1833), .Y(n202) );
  OA222X1_RVT U2152 ( .A1(n2469), .A2(n180), .A3(n181), .A4(n1181), .A5(n2454), 
        .A6(n1833), .Y(n198) );
  OA222X1_RVT U2153 ( .A1(n2468), .A2(n180), .A3(n181), .A4(n1182), .A5(n2453), 
        .A6(n1833), .Y(n194) );
  OA222X1_RVT U2154 ( .A1(n2467), .A2(n180), .A3(n181), .A4(n1183), .A5(n2452), 
        .A6(n1833), .Y(n190) );
  OA222X1_RVT U2155 ( .A1(n2466), .A2(n180), .A3(n181), .A4(n1184), .A5(n2451), 
        .A6(n1833), .Y(n186) );
  OA222X1_RVT U2156 ( .A1(n2464), .A2(n180), .A3(n181), .A4(n1185), .A5(n2446), 
        .A6(n1833), .Y(n178) );
  OR2X1_RVT U2157 ( .A1(n383), .A2(n384), .Y(n175) );
  OR2X1_RVT U2158 ( .A1(n381), .A2(n382), .Y(n169) );
  AO22X1_RVT U2159 ( .A1(n164), .A2(n2474), .A3(n2448), .A4(n239), .Y(n349) );
  AO22X1_RVT U2160 ( .A1(N2243), .A2(n1837), .A3(N2463), .A4(n1463), .Y(n325)
         );
  AO221X1_RVT U2161 ( .A1(N2295), .A2(n1832), .A3(tmp_m1[24]), .A4(n1841), 
        .A5(n327), .Y(n326) );
  AO22X1_RVT U2162 ( .A1(tmp_m1[1]), .A2(n213), .A3(N2515), .A4(n1829), .Y(
        n324) );
  AO22X1_RVT U2163 ( .A1(N2244), .A2(n1837), .A3(N2464), .A4(n1463), .Y(n321)
         );
  AO221X1_RVT U2164 ( .A1(N2296), .A2(n1831), .A3(tmp_m1[25]), .A4(n1840), 
        .A5(n323), .Y(n322) );
  AO22X1_RVT U2165 ( .A1(tmp_m1[2]), .A2(n213), .A3(N2516), .A4(n1828), .Y(
        n320) );
  AO22X1_RVT U2166 ( .A1(N2246), .A2(n1836), .A3(N2466), .A4(n1838), .Y(n313)
         );
  AO221X1_RVT U2167 ( .A1(N2298), .A2(n1832), .A3(tmp_m1[27]), .A4(n1839), 
        .A5(n315), .Y(n314) );
  AO22X1_RVT U2168 ( .A1(tmp_m1[4]), .A2(n213), .A3(N2518), .A4(n1828), .Y(
        n312) );
  AO22X1_RVT U2169 ( .A1(N2250), .A2(n1837), .A3(N2470), .A4(n1463), .Y(n297)
         );
  AO221X1_RVT U2170 ( .A1(N2302), .A2(n1831), .A3(tmp_m1[31]), .A4(n1840), 
        .A5(n299), .Y(n298) );
  AO22X1_RVT U2171 ( .A1(tmp_m1[8]), .A2(n213), .A3(N2522), .A4(n1829), .Y(
        n296) );
  AO22X1_RVT U2172 ( .A1(N2251), .A2(n1837), .A3(N2471), .A4(n1463), .Y(n293)
         );
  AO221X1_RVT U2173 ( .A1(N2303), .A2(n1830), .A3(tmp_m1[32]), .A4(n1841), 
        .A5(n295), .Y(n294) );
  AO22X1_RVT U2174 ( .A1(tmp_m1[9]), .A2(n213), .A3(N2523), .A4(n1827), .Y(
        n292) );
  AO22X1_RVT U2175 ( .A1(N2252), .A2(n1836), .A3(N2472), .A4(n1838), .Y(n289)
         );
  AO221X1_RVT U2176 ( .A1(N2304), .A2(n1831), .A3(tmp_m1[33]), .A4(n1840), 
        .A5(n291), .Y(n290) );
  AO22X1_RVT U2177 ( .A1(tmp_m1[10]), .A2(n213), .A3(N2524), .A4(n1827), .Y(
        n288) );
  AO22X1_RVT U2178 ( .A1(N2253), .A2(n1836), .A3(N2473), .A4(n1838), .Y(n285)
         );
  AO221X1_RVT U2179 ( .A1(N2305), .A2(n1830), .A3(tmp_m1[34]), .A4(n1839), 
        .A5(n287), .Y(n286) );
  AO22X1_RVT U2180 ( .A1(tmp_m1[11]), .A2(n213), .A3(N2525), .A4(n1827), .Y(
        n284) );
  AO22X1_RVT U2181 ( .A1(N2255), .A2(n1836), .A3(N2475), .A4(n1838), .Y(n277)
         );
  AO221X1_RVT U2182 ( .A1(N2307), .A2(n1830), .A3(tmp_m1[36]), .A4(n1839), 
        .A5(n279), .Y(n278) );
  AO22X1_RVT U2183 ( .A1(tmp_m1[13]), .A2(n213), .A3(N2527), .A4(n1827), .Y(
        n276) );
  AO22X1_RVT U2184 ( .A1(N2257), .A2(n1837), .A3(N2477), .A4(n1838), .Y(n269)
         );
  AO221X1_RVT U2185 ( .A1(N2309), .A2(n1832), .A3(tmp_m1[38]), .A4(n1839), 
        .A5(n271), .Y(n270) );
  AO22X1_RVT U2186 ( .A1(tmp_m1[15]), .A2(n213), .A3(N2529), .A4(n1829), .Y(
        n268) );
  AO22X1_RVT U2187 ( .A1(N2258), .A2(n1837), .A3(N2478), .A4(n1838), .Y(n265)
         );
  AO221X1_RVT U2188 ( .A1(N2310), .A2(n1831), .A3(tmp_m1[39]), .A4(n1839), 
        .A5(n267), .Y(n266) );
  AO22X1_RVT U2189 ( .A1(tmp_m1[16]), .A2(n213), .A3(N2530), .A4(n1829), .Y(
        n264) );
  AO22X1_RVT U2190 ( .A1(N2259), .A2(n1837), .A3(N2479), .A4(n1838), .Y(n261)
         );
  AO221X1_RVT U2191 ( .A1(N2311), .A2(n1830), .A3(tmp_m1[40]), .A4(n1840), 
        .A5(n263), .Y(n262) );
  AO22X1_RVT U2192 ( .A1(tmp_m1[17]), .A2(n213), .A3(N2531), .A4(n1828), .Y(
        n260) );
  AO22X1_RVT U2193 ( .A1(N2264), .A2(n1836), .A3(N2484), .A4(n1463), .Y(n230)
         );
  AO221X1_RVT U2194 ( .A1(N2316), .A2(n1831), .A3(tmp_m1[45]), .A4(n1840), 
        .A5(n232), .Y(n231) );
  AO22X1_RVT U2195 ( .A1(N2254), .A2(n1836), .A3(N2474), .A4(n1838), .Y(n281)
         );
  AO221X1_RVT U2196 ( .A1(N2306), .A2(n1832), .A3(tmp_m1[35]), .A4(n1841), 
        .A5(n283), .Y(n282) );
  AO22X1_RVT U2197 ( .A1(tmp_m1[12]), .A2(n1835), .A3(N2526), .A4(n1829), .Y(
        n280) );
  AO22X1_RVT U2198 ( .A1(N2248), .A2(n1836), .A3(N2468), .A4(n1463), .Y(n305)
         );
  AO221X1_RVT U2199 ( .A1(N2300), .A2(n1830), .A3(tmp_m1[29]), .A4(n1840), 
        .A5(n307), .Y(n306) );
  AO22X1_RVT U2200 ( .A1(tmp_m1[6]), .A2(n1835), .A3(N2520), .A4(n1828), .Y(
        n304) );
  AO22X1_RVT U2201 ( .A1(N2262), .A2(n1836), .A3(N2482), .A4(n1463), .Y(n249)
         );
  AO221X1_RVT U2202 ( .A1(N2314), .A2(n1830), .A3(tmp_m1[43]), .A4(n1840), 
        .A5(n251), .Y(n250) );
  AO22X1_RVT U2203 ( .A1(tmp_m1[20]), .A2(n1835), .A3(N2534), .A4(n1829), .Y(
        n248) );
  AO22X1_RVT U2204 ( .A1(N2245), .A2(n1836), .A3(N2465), .A4(n1463), .Y(n317)
         );
  AO221X1_RVT U2205 ( .A1(N2297), .A2(n1832), .A3(tmp_m1[26]), .A4(n1840), 
        .A5(n319), .Y(n318) );
  AO22X1_RVT U2206 ( .A1(tmp_m1[3]), .A2(n1835), .A3(N2517), .A4(n1828), .Y(
        n316) );
  AO22X1_RVT U2207 ( .A1(N2247), .A2(n1837), .A3(N2467), .A4(n1838), .Y(n309)
         );
  AO221X1_RVT U2208 ( .A1(N2299), .A2(n1831), .A3(tmp_m1[28]), .A4(n1839), 
        .A5(n311), .Y(n310) );
  AO22X1_RVT U2209 ( .A1(tmp_m1[5]), .A2(n1835), .A3(N2519), .A4(n1828), .Y(
        n308) );
  AO22X1_RVT U2210 ( .A1(N2249), .A2(n1837), .A3(N2469), .A4(n1463), .Y(n301)
         );
  AO221X1_RVT U2211 ( .A1(N2301), .A2(n1831), .A3(tmp_m1[30]), .A4(n1839), 
        .A5(n303), .Y(n302) );
  AO22X1_RVT U2212 ( .A1(tmp_m1[7]), .A2(n1835), .A3(N2521), .A4(n1827), .Y(
        n300) );
  AO22X1_RVT U2213 ( .A1(N2256), .A2(n1836), .A3(N2476), .A4(n1838), .Y(n273)
         );
  AO221X1_RVT U2214 ( .A1(N2308), .A2(n1830), .A3(tmp_m1[37]), .A4(n1840), 
        .A5(n275), .Y(n274) );
  AO22X1_RVT U2215 ( .A1(tmp_m1[14]), .A2(n1835), .A3(N2528), .A4(n1829), .Y(
        n272) );
  AO22X1_RVT U2216 ( .A1(N2260), .A2(n1837), .A3(N2480), .A4(n1838), .Y(n257)
         );
  AO221X1_RVT U2217 ( .A1(N2312), .A2(n1832), .A3(tmp_m1[41]), .A4(n1839), 
        .A5(n259), .Y(n258) );
  AO22X1_RVT U2218 ( .A1(tmp_m1[18]), .A2(n1835), .A3(N2532), .A4(n1827), .Y(
        n256) );
  AO22X1_RVT U2219 ( .A1(N2261), .A2(n1837), .A3(N2481), .A4(n1463), .Y(n253)
         );
  AO221X1_RVT U2220 ( .A1(N2313), .A2(n1831), .A3(tmp_m1[42]), .A4(n1840), 
        .A5(n255), .Y(n254) );
  AO22X1_RVT U2221 ( .A1(tmp_m1[19]), .A2(n1835), .A3(N2533), .A4(n1828), .Y(
        n252) );
  AO22X1_RVT U2222 ( .A1(N2263), .A2(n1836), .A3(N2483), .A4(n1463), .Y(n245)
         );
  AO22X1_RVT U2223 ( .A1(tmp_m1[21]), .A2(n1835), .A3(N2535), .A4(n1827), .Y(
        n244) );
  OAI22X1_RVT U2224 ( .A1(\sel_2[1] ), .A2(n153), .A3(n154), .A4(n2477), .Y(
        N2800) );
  OA21X1_RVT U2225 ( .A1(n156), .A2(n157), .A3(n158), .Y(n154) );
  OA222X1_RVT U2226 ( .A1(n159), .A2(n2461), .A3(n161), .A4(n2471), .A5(n163), 
        .A6(n2477), .Y(n153) );
  AO21X1_RVT U2227 ( .A1(tmp_m0[24]), .A2(n1560), .A3(n1864), .Y(n619) );
  OR3X2_RVT U2228 ( .A1(n239), .A2(tmp_m1[23]), .A3(n157), .Y(n1782) );
  AO221X1_RVT U2229 ( .A1(tmp_m0[28]), .A2(n620), .A3(tmp_m0[29]), .A4(n619), 
        .A5(n636), .Y(N2093) );
  AO221X1_RVT U2230 ( .A1(n634), .A2(n1851), .A3(tmp_m0[28]), .A4(n617), .A5(
        n635), .Y(N2094) );
  AO22X1_RVT U2231 ( .A1(tmp_m0[30]), .A2(n619), .A3(tmp_m0[29]), .A4(n620), 
        .Y(n635) );
  AO22X1_RVT U2232 ( .A1(tmp_b_m1[7]), .A2(n1952), .A3(n1236), .A4(n1976), .Y(
        n1350) );
  AO22X1_RVT U2233 ( .A1(tmp_b_m1[8]), .A2(n1952), .A3(n1237), .A4(n1976), .Y(
        n1352) );
  AO22X1_RVT U2234 ( .A1(tmp_b_m1[9]), .A2(n1953), .A3(n1238), .A4(n1976), .Y(
        n1354) );
  AO22X1_RVT U2235 ( .A1(tmp_b_m1[10]), .A2(n1953), .A3(n1239), .A4(n1976), 
        .Y(n1356) );
  AO22X1_RVT U2236 ( .A1(tmp_b_m1[11]), .A2(n1953), .A3(n1240), .A4(n1976), 
        .Y(n1358) );
  AO22X1_RVT U2237 ( .A1(tmp_b_m1[12]), .A2(n1953), .A3(n1241), .A4(n1976), 
        .Y(n1360) );
  AO22X1_RVT U2238 ( .A1(tmp_b_m1[13]), .A2(n1953), .A3(n1242), .A4(n1976), 
        .Y(n1362) );
  AO22X1_RVT U2239 ( .A1(tmp_b_m1[14]), .A2(n1953), .A3(n1243), .A4(n1976), 
        .Y(n1364) );
  AO22X1_RVT U2240 ( .A1(tmp_b_m1[15]), .A2(n1953), .A3(n1244), .A4(n1976), 
        .Y(n1366) );
  AO22X1_RVT U2241 ( .A1(tmp_b_m1[16]), .A2(n1953), .A3(n1245), .A4(n1976), 
        .Y(n1368) );
  AO22X1_RVT U2242 ( .A1(tmp_b_m1[17]), .A2(n1953), .A3(n1246), .A4(n1976), 
        .Y(n1370) );
  AO22X1_RVT U2243 ( .A1(tmp_b_m1[18]), .A2(n1953), .A3(n1247), .A4(n1976), 
        .Y(n1372) );
  AO22X1_RVT U2244 ( .A1(tmp_b_m1[19]), .A2(n1953), .A3(n1248), .A4(n1976), 
        .Y(n1374) );
  AO22X1_RVT U2245 ( .A1(tmp_b_m1[20]), .A2(n1953), .A3(n1249), .A4(n1976), 
        .Y(n1376) );
  AO22X1_RVT U2246 ( .A1(tmp_b_m1[21]), .A2(n1953), .A3(n1250), .A4(n1976), 
        .Y(n1378) );
  AO22X1_RVT U2247 ( .A1(tmp_b_m1[22]), .A2(n1954), .A3(n1251), .A4(n1976), 
        .Y(n1380) );
  AO22X1_RVT U2248 ( .A1(tmp_a_e1[0]), .A2(n1954), .A3(n1252), .A4(n1976), .Y(
        n1382) );
  AO22X1_RVT U2249 ( .A1(n1252), .A2(n1954), .A3(a_e[0]), .A4(n1976), .Y(n1383) );
  AO22X1_RVT U2250 ( .A1(tmp_a_e1[1]), .A2(n1954), .A3(n1254), .A4(n1976), .Y(
        n1384) );
  AO22X1_RVT U2251 ( .A1(n1254), .A2(n1954), .A3(a_e[1]), .A4(n1976), .Y(n1385) );
  AO22X1_RVT U2252 ( .A1(tmp_a_e1[2]), .A2(n1954), .A3(n1256), .A4(n1976), .Y(
        n1386) );
  AO22X1_RVT U2253 ( .A1(n1256), .A2(n1954), .A3(a_e[2]), .A4(n1976), .Y(n1387) );
  AO22X1_RVT U2254 ( .A1(tmp_b_e1[3]), .A2(n1949), .A3(n1194), .A4(n1977), .Y(
        n1275) );
  AO22X1_RVT U2255 ( .A1(tmp_b_e1[4]), .A2(n1949), .A3(n1196), .A4(n1977), .Y(
        n1276) );
  AO22X1_RVT U2256 ( .A1(tmp_b_e1[5]), .A2(n1949), .A3(n1198), .A4(n1977), .Y(
        n1277) );
  AO22X1_RVT U2257 ( .A1(tmp_b_e1[6]), .A2(n1949), .A3(n1200), .A4(n1977), .Y(
        n1278) );
  AO22X1_RVT U2258 ( .A1(tmp_b_e1[7]), .A2(n1949), .A3(n1202), .A4(n1977), .Y(
        n1279) );
  AO22X1_RVT U2259 ( .A1(n1188), .A2(n1949), .A3(b_e[0]), .A4(n1977), .Y(n1280) );
  AO22X1_RVT U2260 ( .A1(n1190), .A2(n1949), .A3(b_e[1]), .A4(n1977), .Y(n1281) );
  AO22X1_RVT U2261 ( .A1(n1192), .A2(n1949), .A3(b_e[2]), .A4(n1977), .Y(n1282) );
  AO22X1_RVT U2262 ( .A1(n1194), .A2(n1950), .A3(b_e[3]), .A4(n1977), .Y(n1283) );
  AO22X1_RVT U2263 ( .A1(n1196), .A2(n1950), .A3(b_e[4]), .A4(n1977), .Y(n1284) );
  AO22X1_RVT U2264 ( .A1(n1198), .A2(n1950), .A3(b_e[5]), .A4(n1977), .Y(n1285) );
  AO22X1_RVT U2265 ( .A1(n1200), .A2(n1950), .A3(b_e[6]), .A4(n1977), .Y(n1286) );
  AO22X1_RVT U2266 ( .A1(n1202), .A2(n1950), .A3(b_e[7]), .A4(n1977), .Y(n1287) );
  AO22X1_RVT U2267 ( .A1(tmp_a_m1[0]), .A2(n1950), .A3(n1204), .A4(n1977), .Y(
        n1288) );
  AO22X1_RVT U2268 ( .A1(tmp_a_m1[1]), .A2(n1950), .A3(n1205), .A4(n1977), .Y(
        n1290) );
  AO22X1_RVT U2269 ( .A1(tmp_a_m1[2]), .A2(n1950), .A3(n1206), .A4(n1977), .Y(
        n1292) );
  AO22X1_RVT U2270 ( .A1(tmp_a_m1[3]), .A2(n1950), .A3(n1207), .A4(n1977), .Y(
        n1294) );
  AO22X1_RVT U2271 ( .A1(tmp_a_m1[4]), .A2(n1950), .A3(n1208), .A4(n1977), .Y(
        n1296) );
  AO22X1_RVT U2272 ( .A1(tmp_a_m1[5]), .A2(n1950), .A3(n1209), .A4(n1977), .Y(
        n1298) );
  AO22X1_RVT U2273 ( .A1(tmp_a_m1[6]), .A2(n1950), .A3(n1210), .A4(n1977), .Y(
        n1300) );
  AO22X1_RVT U2274 ( .A1(tmp_a_m1[7]), .A2(n1950), .A3(n1211), .A4(n1977), .Y(
        n1302) );
  AO22X1_RVT U2275 ( .A1(tmp_a_m1[8]), .A2(n1951), .A3(n1212), .A4(n1977), .Y(
        n1304) );
  AO22X1_RVT U2276 ( .A1(n1187), .A2(n1949), .A3(n1609), .A4(n1978), .Y(n1271)
         );
  AO22X1_RVT U2277 ( .A1(n1258), .A2(n1954), .A3(a_e[3]), .A4(n1975), .Y(n1389) );
  AO22X1_RVT U2278 ( .A1(n1260), .A2(n1954), .A3(a_e[4]), .A4(n1975), .Y(n1391) );
  AO22X1_RVT U2279 ( .A1(n1262), .A2(n1954), .A3(a_e[5]), .A4(n1975), .Y(n1393) );
  AO22X1_RVT U2280 ( .A1(n1264), .A2(rst), .A3(a_e[6]), .A4(n1975), .Y(n1395)
         );
  AO22X1_RVT U2281 ( .A1(n1266), .A2(n1949), .A3(a_e[7]), .A4(n1975), .Y(n1397) );
  AO22X1_RVT U2282 ( .A1(n1227), .A2(n1952), .A3(n1605), .A4(n1978), .Y(n1335)
         );
  AO22X1_RVT U2283 ( .A1(sel_1[0]), .A2(n1978), .A3(n1186), .A4(n1948), .Y(
        n1268) );
  AO22X1_RVT U2284 ( .A1(\sel_2[1] ), .A2(n1948), .A3(sel_1[1]), .A4(n1978), 
        .Y(n1269) );
  AO22X1_RVT U2285 ( .A1(tmp_b_s1), .A2(n1948), .A3(n1187), .A4(n1978), .Y(
        n1270) );
  AO22X1_RVT U2286 ( .A1(tmp_a_e1[7]), .A2(n1948), .A3(n1266), .A4(n1975), .Y(
        n1396) );
  AO22X1_RVT U2287 ( .A1(tmp_b_e1[0]), .A2(n1949), .A3(n1188), .A4(n1978), .Y(
        n1272) );
  AO22X1_RVT U2288 ( .A1(tmp_b_e1[1]), .A2(n1949), .A3(n1190), .A4(n1978), .Y(
        n1273) );
  AO22X1_RVT U2289 ( .A1(tmp_b_e1[2]), .A2(n1949), .A3(n1192), .A4(n1978), .Y(
        n1274) );
  AO22X1_RVT U2290 ( .A1(tmp_a_m1[9]), .A2(n1951), .A3(n1213), .A4(n1978), .Y(
        n1306) );
  AO22X1_RVT U2291 ( .A1(tmp_a_m1[10]), .A2(n1951), .A3(n1214), .A4(n1955), 
        .Y(n1308) );
  AO22X1_RVT U2292 ( .A1(tmp_a_m1[11]), .A2(n1951), .A3(n1215), .A4(n1978), 
        .Y(n1310) );
  AO22X1_RVT U2293 ( .A1(tmp_a_m1[12]), .A2(n1951), .A3(n1216), .A4(n1955), 
        .Y(n1312) );
  AO22X1_RVT U2294 ( .A1(tmp_a_m1[13]), .A2(n1951), .A3(n1217), .A4(n1975), 
        .Y(n1314) );
  AO22X1_RVT U2295 ( .A1(tmp_a_m1[14]), .A2(n1951), .A3(n1218), .A4(n1978), 
        .Y(n1316) );
  AO22X1_RVT U2296 ( .A1(tmp_a_m1[15]), .A2(n1951), .A3(n1219), .A4(n1955), 
        .Y(n1318) );
  AO22X1_RVT U2297 ( .A1(tmp_a_m1[16]), .A2(n1951), .A3(n1220), .A4(n1978), 
        .Y(n1320) );
  AO22X1_RVT U2298 ( .A1(tmp_a_m1[17]), .A2(n1951), .A3(n1221), .A4(n1956), 
        .Y(n1322) );
  AO22X1_RVT U2299 ( .A1(tmp_a_m1[18]), .A2(n1951), .A3(n1222), .A4(n1955), 
        .Y(n1324) );
  AO22X1_RVT U2300 ( .A1(tmp_a_m1[19]), .A2(n1951), .A3(n1223), .A4(n1978), 
        .Y(n1326) );
  AO22X1_RVT U2301 ( .A1(tmp_a_m1[20]), .A2(n1951), .A3(n1224), .A4(n1956), 
        .Y(n1328) );
  AO22X1_RVT U2302 ( .A1(tmp_a_m1[21]), .A2(n1952), .A3(n1225), .A4(n1955), 
        .Y(n1330) );
  AO22X1_RVT U2303 ( .A1(tmp_a_m1[22]), .A2(n1952), .A3(n1226), .A4(n1978), 
        .Y(n1332) );
  AO22X1_RVT U2304 ( .A1(tmp_a_s1), .A2(n1952), .A3(n1227), .A4(n1956), .Y(
        n1334) );
  AO22X1_RVT U2305 ( .A1(tmp_b_m1[0]), .A2(n1952), .A3(n1229), .A4(n1955), .Y(
        n1336) );
  AO22X1_RVT U2306 ( .A1(tmp_b_m1[1]), .A2(n1952), .A3(n1230), .A4(n1978), .Y(
        n1338) );
  AO22X1_RVT U2307 ( .A1(tmp_b_m1[2]), .A2(n1952), .A3(n1231), .A4(n1956), .Y(
        n1340) );
  AO22X1_RVT U2308 ( .A1(tmp_b_m1[3]), .A2(n1952), .A3(n1232), .A4(n1955), .Y(
        n1342) );
  AO22X1_RVT U2309 ( .A1(tmp_b_m1[4]), .A2(n1952), .A3(n1233), .A4(n1978), .Y(
        n1344) );
  AO22X1_RVT U2310 ( .A1(tmp_b_m1[5]), .A2(n1952), .A3(n1234), .A4(n1956), .Y(
        n1346) );
  AO22X1_RVT U2311 ( .A1(tmp_b_m1[6]), .A2(n1952), .A3(n1235), .A4(n1955), .Y(
        n1348) );
  AO22X1_RVT U2312 ( .A1(tmp_a_e1[3]), .A2(n1954), .A3(n1258), .A4(n1975), .Y(
        n1388) );
  AO22X1_RVT U2313 ( .A1(tmp_a_e1[4]), .A2(n1954), .A3(n1260), .A4(n1975), .Y(
        n1390) );
  AO22X1_RVT U2314 ( .A1(tmp_a_e1[5]), .A2(n1954), .A3(n1262), .A4(n1975), .Y(
        n1392) );
  AO22X1_RVT U2315 ( .A1(n1854), .A2(tmp_b_m1[1]), .A3(n1558), .A4(tmp_a_m1[1]), .Y(n327) );
  AO22X1_RVT U2316 ( .A1(n1854), .A2(tmp_b_m1[2]), .A3(n1558), .A4(tmp_a_m1[2]), .Y(n323) );
  AO22X1_RVT U2317 ( .A1(n1854), .A2(tmp_b_m1[3]), .A3(n1558), .A4(tmp_a_m1[3]), .Y(n319) );
  AO22X1_RVT U2318 ( .A1(n1854), .A2(tmp_b_m1[4]), .A3(n1558), .A4(tmp_a_m1[4]), .Y(n315) );
  AO22X1_RVT U2319 ( .A1(n1854), .A2(tmp_b_m1[5]), .A3(n1558), .A4(tmp_a_m1[5]), .Y(n311) );
  AO22X1_RVT U2320 ( .A1(n1854), .A2(tmp_b_m1[6]), .A3(n1558), .A4(tmp_a_m1[6]), .Y(n307) );
  AO22X1_RVT U2321 ( .A1(n1854), .A2(tmp_b_m1[7]), .A3(n1558), .A4(tmp_a_m1[7]), .Y(n303) );
  AO22X1_RVT U2322 ( .A1(n1854), .A2(tmp_b_m1[8]), .A3(n1558), .A4(tmp_a_m1[8]), .Y(n299) );
  AO22X1_RVT U2323 ( .A1(n1854), .A2(tmp_b_m1[9]), .A3(n1558), .A4(tmp_a_m1[9]), .Y(n295) );
  AO22X1_RVT U2324 ( .A1(n1854), .A2(tmp_b_m1[10]), .A3(n1558), .A4(
        tmp_a_m1[10]), .Y(n291) );
  AO22X1_RVT U2325 ( .A1(n1854), .A2(tmp_b_m1[11]), .A3(n1558), .A4(
        tmp_a_m1[11]), .Y(n287) );
  AO22X1_RVT U2326 ( .A1(tmp_a_e1[6]), .A2(rst), .A3(n1264), .A4(n1975), .Y(
        n1394) );
  AO22X1_RVT U2327 ( .A1(n1854), .A2(tmp_b_m1[0]), .A3(n1558), .A4(tmp_a_m1[0]), .Y(N2769) );
  AO22X1_RVT U2328 ( .A1(n1855), .A2(tmp_b_m1[17]), .A3(n1558), .A4(
        tmp_a_m1[17]), .Y(n263) );
  AO22X1_RVT U2329 ( .A1(n1855), .A2(tmp_b_m1[22]), .A3(n1558), .A4(
        tmp_a_m1[22]), .Y(n232) );
  AO22X1_RVT U2330 ( .A1(n1855), .A2(tmp_b_m1[21]), .A3(n1558), .A4(
        tmp_a_m1[21]), .Y(n247) );
  AO22X1_RVT U2331 ( .A1(n1855), .A2(tmp_b_m1[14]), .A3(n1558), .A4(
        tmp_a_m1[14]), .Y(n275) );
  AO22X1_RVT U2332 ( .A1(n1855), .A2(tmp_b_m1[13]), .A3(n1558), .A4(
        tmp_a_m1[13]), .Y(n279) );
  AO22X1_RVT U2333 ( .A1(n1855), .A2(tmp_b_m1[19]), .A3(n1558), .A4(
        tmp_a_m1[19]), .Y(n255) );
  AO22X1_RVT U2334 ( .A1(n1855), .A2(tmp_b_m1[12]), .A3(n1558), .A4(
        tmp_a_m1[12]), .Y(n283) );
  AO22X1_RVT U2335 ( .A1(n1855), .A2(tmp_b_m1[16]), .A3(n1558), .A4(
        tmp_a_m1[16]), .Y(n267) );
  AO22X1_RVT U2336 ( .A1(n1855), .A2(tmp_b_m1[15]), .A3(n1558), .A4(
        tmp_a_m1[15]), .Y(n271) );
  AO22X1_RVT U2337 ( .A1(n1855), .A2(tmp_b_m1[18]), .A3(n1558), .A4(
        tmp_a_m1[18]), .Y(n259) );
  AO22X1_RVT U2338 ( .A1(n1855), .A2(tmp_b_m1[20]), .A3(n1558), .A4(
        tmp_a_m1[20]), .Y(n251) );
  OA21X1_RVT U2339 ( .A1(tmp_e1[8]), .A2(n1783), .A3(n1784), .Y(N2233) );
  AND4X1_RVT U2340 ( .A1(tmp_e1[1]), .A2(tmp_e1[5]), .A3(tmp_e1[2]), .A4(n2421), .Y(n1783) );
  INVX1_RVT U2341 ( .A(rst), .Y(n1956) );
  INVX1_RVT U2342 ( .A(rst), .Y(n1955) );
  AO221X1_RVT U2343 ( .A1(N2315), .A2(n1830), .A3(tmp_m1[44]), .A4(n1839), 
        .A5(n247), .Y(n246) );
  INVX1_RVT U2344 ( .A(n1834), .Y(n1835) );
  INVX1_RVT U2345 ( .A(n213), .Y(n1834) );
  NBUFFX2_RVT U2346 ( .A(n2319), .Y(n1812) );
  NAND2X0_RVT U2347 ( .A1(n1593), .A2(tmp_m0[3]), .Y(n428) );
  AO222X1_RVT U2348 ( .A1(n1912), .A2(n2480), .A3(n1912), .A4(n2482), .A5(
        N1129), .A6(n1765), .Y(n990) );
  OA222X1_RVT U2349 ( .A1(n1894), .A2(n1787), .A3(n648), .A4(n1788), .A5(n1861), .A6(n1789), .Y(n561) );
  AND4X1_RVT U2350 ( .A1(n563), .A2(n564), .A3(n565), .A4(n566), .Y(n1788) );
  OA22X1_RVT U2351 ( .A1(n1504), .A2(n1822), .A3(n1690), .A4(n1819), .Y(n564)
         );
  AO221X1_RVT U2352 ( .A1(n556), .A2(n1850), .A3(tmp_m0[39]), .A4(n1857), .A5(
        n557), .Y(N2104) );
  OA222X1_RVT U2353 ( .A1(n1795), .A2(n1861), .A3(n1794), .A4(n1604), .A5(n648), .A6(n1796), .Y(n392) );
  AND4X1_RVT U2354 ( .A1(n398), .A2(n399), .A3(n400), .A4(n401), .Y(n1796) );
  OA22X1_RVT U2355 ( .A1(n426), .A2(n2316), .A3(n428), .A4(n1475), .Y(n420) );
  OR2X1_RVT U2356 ( .A1(n2149), .A2(tmp_m0[2]), .Y(n432) );
  INVX1_RVT U2357 ( .A(n2290), .Y(n2124) );
  OR2X1_RVT U2358 ( .A1(n648), .A2(n408), .Y(n577) );
  NAND2X0_RVT U2359 ( .A1(tmp_m0[11]), .A2(n1519), .Y(n408) );
  INVX1_RVT U2360 ( .A(tmp_m0[11]), .Y(n2300) );
  INVX1_RVT U2361 ( .A(tmp_m0[9]), .Y(n2302) );
  INVX1_RVT U2362 ( .A(tmp_m0[7]), .Y(n2296) );
  INVX1_RVT U2363 ( .A(tmp_m0[26]), .Y(n2132) );
  INVX1_RVT U2364 ( .A(tmp_m0[1]), .Y(n2289) );
  INVX1_RVT U2365 ( .A(tmp_m0[2]), .Y(n2287) );
  INVX1_RVT U2366 ( .A(tmp_m0[3]), .Y(n2291) );
  INVX0_RVT U2367 ( .A(sel_0[0]), .Y(n2325) );
  NAND2X0_RVT U2368 ( .A1(sel_0[1]), .A2(n2325), .Y(n1153) );
  NAND2X0_RVT U2369 ( .A1(n1153), .A2(sel_0[1]), .Y(n1154) );
  NAND2X0_RVT U2370 ( .A1(n1490), .A2(n1573), .Y(n1981) );
  OA21X1_RVT U2371 ( .A1(b_m[1]), .A2(n1582), .A3(n1928), .Y(n1979) );
  AO22X1_RVT U2372 ( .A1(b_m[1]), .A2(n1582), .A3(n1979), .A4(n1517), .Y(n1980) );
  AO222X1_RVT U2373 ( .A1(n1930), .A2(n1581), .A3(n1981), .A4(n1980), .A5(
        b_m[3]), .A6(n1562), .Y(n1982) );
  OA221X1_RVT U2374 ( .A1(b_m[3]), .A2(n1562), .A3(b_m[4]), .A4(n1576), .A5(
        n1982), .Y(n1983) );
  AO221X1_RVT U2375 ( .A1(b_m[4]), .A2(n1576), .A3(n1931), .A4(n1563), .A5(
        n1983), .Y(n1984) );
  OA221X1_RVT U2376 ( .A1(n1931), .A2(n1563), .A3(b_m[6]), .A4(n1577), .A5(
        n1984), .Y(n1985) );
  AO221X1_RVT U2377 ( .A1(b_m[6]), .A2(n1577), .A3(b_m[7]), .A4(n1564), .A5(
        n1985), .Y(n1986) );
  OA221X1_RVT U2378 ( .A1(b_m[7]), .A2(n1564), .A3(n1932), .A4(n1578), .A5(
        n1986), .Y(n1987) );
  AO221X1_RVT U2379 ( .A1(n1932), .A2(n1578), .A3(b_m[9]), .A4(n1513), .A5(
        n1987), .Y(n1988) );
  OA221X1_RVT U2380 ( .A1(b_m[9]), .A2(n1513), .A3(b_m[10]), .A4(n1580), .A5(
        n1988), .Y(n1989) );
  AO221X1_RVT U2381 ( .A1(b_m[10]), .A2(n1580), .A3(b_m[11]), .A4(n1514), .A5(
        n1989), .Y(n1990) );
  OA221X1_RVT U2382 ( .A1(b_m[11]), .A2(n1514), .A3(b_m[12]), .A4(n1575), .A5(
        n1990), .Y(n1991) );
  AO221X1_RVT U2383 ( .A1(b_m[12]), .A2(n1575), .A3(n1410), .A4(n1569), .A5(
        n1991), .Y(n1992) );
  OA221X1_RVT U2384 ( .A1(n1410), .A2(n1569), .A3(b_m[14]), .A4(n1570), .A5(
        n1992), .Y(n1993) );
  AO221X1_RVT U2385 ( .A1(b_m[14]), .A2(n1570), .A3(b_m[15]), .A4(n1565), .A5(
        n1993), .Y(n1994) );
  OA221X1_RVT U2386 ( .A1(b_m[15]), .A2(n1565), .A3(n1934), .A4(n1579), .A5(
        n1994), .Y(n1995) );
  AO221X1_RVT U2387 ( .A1(n1934), .A2(n1579), .A3(n1936), .A4(n1566), .A5(
        n1995), .Y(n1996) );
  OA221X1_RVT U2388 ( .A1(n1936), .A2(n1566), .A3(b_m[18]), .A4(n1571), .A5(
        n1996), .Y(n1997) );
  AO221X1_RVT U2389 ( .A1(b_m[18]), .A2(n1571), .A3(b_m[19]), .A4(n1567), .A5(
        n1997), .Y(n1998) );
  OA221X1_RVT U2390 ( .A1(b_m[19]), .A2(n1567), .A3(b_m[20]), .A4(n1512), .A5(
        n1998), .Y(n1999) );
  AO221X1_RVT U2391 ( .A1(b_m[20]), .A2(n1512), .A3(n1938), .A4(n1568), .A5(
        n1999), .Y(n2000) );
  OA221X1_RVT U2392 ( .A1(n1938), .A2(n1568), .A3(b_m[22]), .A4(n1572), .A5(
        n2000), .Y(n2001) );
  AO21X1_RVT U2393 ( .A1(b_m[22]), .A2(n1572), .A3(n2001), .Y(n2003) );
  NAND2X0_RVT U2394 ( .A1(a_m[23]), .A2(n1574), .Y(n2002) );
  AO22X1_RVT U2395 ( .A1(n1467), .A2(n1515), .A3(n2003), .A4(n2002), .Y(n2004)
         );
  NAND3X0_RVT U2396 ( .A1(n2436), .A2(n2439), .A3(n2004), .Y(n1176) );
  NAND2X0_RVT U2397 ( .A1(n2324), .A2(n1147), .Y(n1140) );
  NAND2X0_RVT U2398 ( .A1(n2016), .A2(n1147), .Y(n1143) );
  AO22X1_RVT U2399 ( .A1(n2440), .A2(N374), .A3(N458), .A4(n2323), .Y(n2008)
         );
  INVX0_RVT U2400 ( .A(n1147), .Y(n2326) );
  AO22X1_RVT U2401 ( .A1(N94), .A2(N374), .A3(N458), .A4(n2324), .Y(n2007) );
  AO22X1_RVT U2402 ( .A1(n2005), .A2(n2325), .A3(n1781), .A4(n2016), .Y(n2012)
         );
  AO22X1_RVT U2403 ( .A1(n1031), .A2(n2325), .A3(n2438), .A4(n1781), .Y(n2015)
         );
  AO22X1_RVT U2404 ( .A1(N483), .A2(n2012), .A3(N432), .A4(n2015), .Y(n2006)
         );
  AO221X1_RVT U2405 ( .A1(n2008), .A2(n2325), .A3(n1781), .A4(n2007), .A5(
        n2006), .Y(n2009) );
  NAND2X0_RVT U2406 ( .A1(n2009), .A2(n1516), .Y(n2010) );
  NAND2X0_RVT U2407 ( .A1(n2323), .A2(n2325), .Y(n2013) );
  AOI21X1_RVT U2408 ( .A1(n1141), .A2(n2013), .A3(sel_0[1]), .Y(net27435) );
  NAND2X0_RVT U2409 ( .A1(n2015), .A2(n1516), .Y(net27586) );
  AND2X1_RVT U2410 ( .A1(n2438), .A2(n2326), .Y(n2019) );
  MUX21X1_RVT U2411 ( .A1(n2019), .A2(n1031), .S0(sel_0[0]), .Y(n2020) );
  NAND2X0_RVT U2412 ( .A1(n2020), .A2(n1516), .Y(net27580) );
  AO22X1_RVT U2413 ( .A1(N1010), .A2(net32880), .A3(N953), .A4(net32864), .Y(
        n2021) );
  AO22X1_RVT U2414 ( .A1(N165), .A2(net32924), .A3(N474), .A4(net32956), .Y(
        n2025) );
  AO222X1_RVT U2415 ( .A1(N449), .A2(net27435), .A3(N365), .A4(net32950), .A5(
        N423), .A6(net32962), .Y(n2024) );
  AO22X1_RVT U2416 ( .A1(N1009), .A2(net32882), .A3(N952), .A4(net32870), .Y(
        n2022) );
  AO221X1_RVT U2417 ( .A1(N249), .A2(net32930), .A3(N223), .A4(net32938), .A5(
        n2022), .Y(n2023) );
  OR3X1_RVT U2418 ( .A1(n2025), .A2(n2024), .A3(n2023), .Y(N1067) );
  AO22X1_RVT U2419 ( .A1(N1007), .A2(net32882), .A3(N950), .A4(net32870), .Y(
        n2026) );
  AO221X1_RVT U2420 ( .A1(N247), .A2(net32930), .A3(N221), .A4(net27434), .A5(
        n2026), .Y(n2027) );
  AO22X1_RVT U2421 ( .A1(N164), .A2(net32924), .A3(N473), .A4(net32956), .Y(
        n2031) );
  AO222X1_RVT U2422 ( .A1(N448), .A2(net27435), .A3(N364), .A4(net32950), .A5(
        N422), .A6(net32962), .Y(n2030) );
  AO22X1_RVT U2423 ( .A1(N1008), .A2(net32882), .A3(N951), .A4(net32870), .Y(
        n2028) );
  OR3X1_RVT U2424 ( .A1(n2031), .A2(n2030), .A3(n2029), .Y(N1066) );
  AO22X1_RVT U2425 ( .A1(N162), .A2(net32924), .A3(N471), .A4(net32956), .Y(
        n2035) );
  AO222X1_RVT U2426 ( .A1(N446), .A2(net27435), .A3(N362), .A4(net32950), .A5(
        N420), .A6(net32962), .Y(n2034) );
  AO22X1_RVT U2427 ( .A1(N1006), .A2(net32882), .A3(N949), .A4(net32870), .Y(
        n2032) );
  AO221X1_RVT U2428 ( .A1(N246), .A2(net32930), .A3(N220), .A4(net27434), .A5(
        n2032), .Y(n2033) );
  OR3X1_RVT U2429 ( .A1(n2035), .A2(n2034), .A3(n2033), .Y(N1064) );
  AO22X1_RVT U2430 ( .A1(N160), .A2(net32924), .A3(N469), .A4(net32956), .Y(
        n2039) );
  AO222X1_RVT U2431 ( .A1(N444), .A2(net27435), .A3(N360), .A4(net32950), .A5(
        N418), .A6(net32962), .Y(n2038) );
  AO22X1_RVT U2432 ( .A1(N1004), .A2(net32882), .A3(N947), .A4(net32868), .Y(
        n2036) );
  AO221X1_RVT U2433 ( .A1(N244), .A2(net32930), .A3(N218), .A4(net27434), .A5(
        n2036), .Y(n2037) );
  OR3X1_RVT U2434 ( .A1(n2039), .A2(n2038), .A3(n2037), .Y(N1062) );
  AO22X1_RVT U2435 ( .A1(N161), .A2(net32924), .A3(N470), .A4(net32956), .Y(
        n2043) );
  AO222X1_RVT U2436 ( .A1(N445), .A2(net27435), .A3(N361), .A4(net32950), .A5(
        N419), .A6(net32962), .Y(n2042) );
  AO22X1_RVT U2437 ( .A1(N1005), .A2(net32882), .A3(N948), .A4(net32864), .Y(
        n2040) );
  AO221X1_RVT U2438 ( .A1(N245), .A2(net32930), .A3(N219), .A4(net27434), .A5(
        n2040), .Y(n2041) );
  OR3X1_RVT U2439 ( .A1(n2043), .A2(n2042), .A3(n2041), .Y(N1063) );
  NAND3X0_RVT U2440 ( .A1(n1775), .A2(n1613), .A3(n1790), .Y(n2103) );
  AO22X1_RVT U2441 ( .A1(N173), .A2(net32924), .A3(N482), .A4(net32956), .Y(
        n2047) );
  AO222X1_RVT U2442 ( .A1(N457), .A2(net27435), .A3(N373), .A4(net32950), .A5(
        N431), .A6(net32962), .Y(n2046) );
  AO22X1_RVT U2443 ( .A1(N1017), .A2(net32882), .A3(N960), .A4(net32864), .Y(
        n2044) );
  AO221X1_RVT U2444 ( .A1(N257), .A2(net32930), .A3(N231), .A4(net27434), .A5(
        n2044), .Y(n2045) );
  AO222X1_RVT U2445 ( .A1(N961), .A2(net32870), .A3(N232), .A4(net27434), .A5(
        N1018), .A6(net32876), .Y(n2049) );
  AO221X1_RVT U2446 ( .A1(N174), .A2(net32924), .A3(N258), .A4(net32930), .A5(
        n1856), .Y(n2048) );
  OR2X1_RVT U2447 ( .A1(n2049), .A2(n2048), .Y(N1076) );
  AO22X1_RVT U2448 ( .A1(N171), .A2(net32924), .A3(N480), .A4(net32956), .Y(
        n2053) );
  AO222X1_RVT U2449 ( .A1(N455), .A2(net27435), .A3(N371), .A4(net32950), .A5(
        N429), .A6(net32962), .Y(n2052) );
  AO22X1_RVT U2450 ( .A1(N1015), .A2(net32882), .A3(N958), .A4(net32864), .Y(
        n2050) );
  AO221X1_RVT U2451 ( .A1(N255), .A2(net32930), .A3(N229), .A4(net27434), .A5(
        n2050), .Y(n2051) );
  OR3X1_RVT U2452 ( .A1(n2053), .A2(n2052), .A3(n2051), .Y(N1073) );
  AO22X1_RVT U2453 ( .A1(N172), .A2(net32924), .A3(N481), .A4(net32956), .Y(
        n2057) );
  AO222X1_RVT U2454 ( .A1(N456), .A2(net27435), .A3(N372), .A4(net32950), .A5(
        N430), .A6(net32962), .Y(n2056) );
  AO22X1_RVT U2455 ( .A1(N1016), .A2(net32882), .A3(N959), .A4(net32864), .Y(
        n2054) );
  AO221X1_RVT U2456 ( .A1(N256), .A2(net32930), .A3(N230), .A4(net27434), .A5(
        n2054), .Y(n2055) );
  OR3X1_RVT U2457 ( .A1(n2057), .A2(n2056), .A3(n2055), .Y(N1074) );
  AO22X1_RVT U2458 ( .A1(N170), .A2(net32924), .A3(N479), .A4(net32956), .Y(
        n2061) );
  AO222X1_RVT U2459 ( .A1(N454), .A2(net32946), .A3(N370), .A4(net32950), .A5(
        N428), .A6(net32962), .Y(n2060) );
  AO22X1_RVT U2460 ( .A1(N1014), .A2(net32882), .A3(N957), .A4(net32864), .Y(
        n2058) );
  AO221X1_RVT U2461 ( .A1(N254), .A2(net32930), .A3(N228), .A4(net27434), .A5(
        n2058), .Y(n2059) );
  OR3X1_RVT U2462 ( .A1(n2061), .A2(n2060), .A3(n2059), .Y(N1072) );
  AO22X1_RVT U2463 ( .A1(N167), .A2(net32926), .A3(N476), .A4(net32956), .Y(
        n2065) );
  AO222X1_RVT U2464 ( .A1(N451), .A2(net27435), .A3(N367), .A4(net32950), .A5(
        N425), .A6(net32962), .Y(n2064) );
  AO22X1_RVT U2465 ( .A1(N1011), .A2(net32882), .A3(N954), .A4(net32864), .Y(
        n2062) );
  AO221X1_RVT U2466 ( .A1(N251), .A2(net32932), .A3(N225), .A4(net27434), .A5(
        n2062), .Y(n2063) );
  OR3X1_RVT U2467 ( .A1(n2065), .A2(n2064), .A3(n2063), .Y(N1069) );
  AO22X1_RVT U2468 ( .A1(N168), .A2(net32926), .A3(N477), .A4(net32958), .Y(
        n2069) );
  AO222X1_RVT U2469 ( .A1(N452), .A2(net32946), .A3(N368), .A4(net32952), .A5(
        N426), .A6(net27438), .Y(n2068) );
  AO22X1_RVT U2470 ( .A1(N1012), .A2(net32882), .A3(N955), .A4(net32864), .Y(
        n2066) );
  AO221X1_RVT U2471 ( .A1(N252), .A2(net32932), .A3(N226), .A4(net32938), .A5(
        n2066), .Y(n2067) );
  OR3X1_RVT U2472 ( .A1(n2069), .A2(n2068), .A3(n2067), .Y(N1070) );
  AO22X1_RVT U2473 ( .A1(N169), .A2(net32926), .A3(N478), .A4(net32958), .Y(
        n2073) );
  AO222X1_RVT U2474 ( .A1(N453), .A2(net32946), .A3(N369), .A4(net32952), .A5(
        N427), .A6(net27438), .Y(n2072) );
  AO22X1_RVT U2475 ( .A1(N1013), .A2(net32882), .A3(N956), .A4(net32864), .Y(
        n2070) );
  AO221X1_RVT U2476 ( .A1(N253), .A2(net32932), .A3(N227), .A4(net32938), .A5(
        n2070), .Y(n2071) );
  OR3X1_RVT U2477 ( .A1(n2073), .A2(n2072), .A3(n2071), .Y(N1071) );
  AO22X1_RVT U2478 ( .A1(N159), .A2(net32926), .A3(N468), .A4(net32958), .Y(
        n2077) );
  AO222X1_RVT U2479 ( .A1(N443), .A2(net32946), .A3(N359), .A4(net32952), .A5(
        net27438), .A6(N417), .Y(n2076) );
  AO22X1_RVT U2480 ( .A1(N1003), .A2(net32880), .A3(N946), .A4(net32864), .Y(
        n2074) );
  AO221X1_RVT U2481 ( .A1(N243), .A2(net32932), .A3(N217), .A4(net32938), .A5(
        n2074), .Y(n2075) );
  OR3X1_RVT U2482 ( .A1(n2077), .A2(n2076), .A3(n2075), .Y(N1061) );
  NAND2X0_RVT U2483 ( .A1(n1585), .A2(n1844), .Y(n2078) );
  NAND3X0_RVT U2484 ( .A1(n1699), .A2(n1493), .A3(n1474), .Y(n2090) );
  NAND4X0_RVT U2485 ( .A1(n1586), .A2(n1468), .A3(n1484), .A4(n1492), .Y(n2089) );
  NAND3X0_RVT U2486 ( .A1(n2088), .A2(n1491), .A3(n1803), .Y(n994) );
  AO22X1_RVT U2487 ( .A1(N157), .A2(net32926), .A3(N466), .A4(net32958), .Y(
        n2082) );
  AO222X1_RVT U2488 ( .A1(N441), .A2(net32946), .A3(N357), .A4(net32952), .A5(
        N415), .A6(net32962), .Y(n2081) );
  AO22X1_RVT U2489 ( .A1(N1001), .A2(net32880), .A3(N944), .A4(net32864), .Y(
        n2079) );
  AO221X1_RVT U2490 ( .A1(N241), .A2(net32932), .A3(N215), .A4(net32938), .A5(
        n2079), .Y(n2080) );
  OR3X1_RVT U2491 ( .A1(n2082), .A2(n2081), .A3(n2080), .Y(N1059) );
  AO22X1_RVT U2492 ( .A1(N158), .A2(net32926), .A3(N467), .A4(net32958), .Y(
        n2086) );
  AO222X1_RVT U2493 ( .A1(N442), .A2(net32946), .A3(N358), .A4(net32952), .A5(
        N416), .A6(net32962), .Y(n2085) );
  AO22X1_RVT U2494 ( .A1(N1002), .A2(net32880), .A3(N945), .A4(net32864), .Y(
        n2083) );
  AO221X1_RVT U2495 ( .A1(N242), .A2(net32932), .A3(N216), .A4(net32938), .A5(
        n2083), .Y(n2084) );
  NAND2X0_RVT U2496 ( .A1(tmp_m0[7]), .A2(n2301), .Y(n2295) );
  NAND2X0_RVT U2497 ( .A1(tmp_m0[8]), .A2(n2322), .Y(n515) );
  NAND3X0_RVT U2498 ( .A1(n1586), .A2(n1492), .A3(n2089), .Y(n647) );
  AO22X1_RVT U2499 ( .A1(N156), .A2(net32926), .A3(N465), .A4(net32958), .Y(
        n2094) );
  AO22X1_RVT U2500 ( .A1(N1000), .A2(net32880), .A3(N943), .A4(net32864), .Y(
        n2092) );
  AO221X1_RVT U2501 ( .A1(N240), .A2(net32932), .A3(N214), .A4(net32938), .A5(
        n2092), .Y(n2093) );
  OR3X1_RVT U2502 ( .A1(n2094), .A2(n1541), .A3(n2093), .Y(N1058) );
  NAND2X0_RVT U2503 ( .A1(tmp_m0[6]), .A2(n1768), .Y(n2293) );
  NAND2X0_RVT U2504 ( .A1(n2095), .A2(n2322), .Y(n486) );
  INVX0_RVT U2505 ( .A(sel_1[1]), .Y(n2318) );
  NAND3X0_RVT U2506 ( .A1(tmp_m0[23]), .A2(sel_1[1]), .A3(n454), .Y(n455) );
  AO221X1_RVT U2507 ( .A1(N965), .A2(net32868), .A3(N1022), .A4(net32876), 
        .A5(n1856), .Y(N1080) );
  AO221X1_RVT U2508 ( .A1(N966), .A2(net32868), .A3(N1023), .A4(net32876), 
        .A5(n1856), .Y(N1081) );
  AO221X1_RVT U2509 ( .A1(N963), .A2(net32868), .A3(N1020), .A4(net32878), 
        .A5(n1856), .Y(N1078) );
  AO221X1_RVT U2510 ( .A1(N964), .A2(net32866), .A3(N1021), .A4(net32878), 
        .A5(n1856), .Y(N1079) );
  AO21X1_RVT U2511 ( .A1(n1878), .A2(n1560), .A3(n1847), .Y(n617) );
  NAND2X0_RVT U2512 ( .A1(n1890), .A2(n1560), .Y(n2139) );
  NAND2X0_RVT U2513 ( .A1(n617), .A2(tmp_m0[27]), .Y(n2097) );
  NAND3X0_RVT U2514 ( .A1(n1851), .A2(n1863), .A3(tmp_m0[25]), .Y(n2096) );
  NAND3X0_RVT U2515 ( .A1(n2098), .A2(n2097), .A3(n2096), .Y(n636) );
  AO221X1_RVT U2516 ( .A1(N967), .A2(net32868), .A3(N1024), .A4(net32878), 
        .A5(n1856), .Y(N1082) );
  AO222X1_RVT U2517 ( .A1(n1890), .A2(tmp_m0[27]), .A3(tmp_m0[26]), .A4(n1863), 
        .A5(tmp_m0[25]), .A6(n1899), .Y(n634) );
  AO221X1_RVT U2518 ( .A1(N968), .A2(net32866), .A3(N1025), .A4(net32878), 
        .A5(n1856), .Y(N1083) );
  AO22X1_RVT U2519 ( .A1(tmp_m0[26]), .A2(n1900), .A3(n1890), .A4(tmp_m0[28]), 
        .Y(n2100) );
  AO221X1_RVT U2520 ( .A1(n1863), .A2(tmp_m0[27]), .A3(tmp_m0[25]), .A4(n1871), 
        .A5(n2100), .Y(n629) );
  AO221X1_RVT U2521 ( .A1(N969), .A2(net32866), .A3(N1026), .A4(net32878), 
        .A5(n1856), .Y(N1084) );
  AO221X1_RVT U2522 ( .A1(N970), .A2(net32866), .A3(N1027), .A4(net32878), 
        .A5(n1856), .Y(N1085) );
  AO221X1_RVT U2523 ( .A1(N971), .A2(net32866), .A3(N1028), .A4(net32878), 
        .A5(n1856), .Y(N1086) );
  AO221X1_RVT U2524 ( .A1(N972), .A2(net32866), .A3(N1029), .A4(net32878), 
        .A5(n1856), .Y(N1087) );
  AO221X1_RVT U2525 ( .A1(N973), .A2(net32866), .A3(N1030), .A4(net32878), 
        .A5(n1856), .Y(N1088) );
  NAND2X0_RVT U2526 ( .A1(n2320), .A2(n2101), .Y(n581) );
  NAND2X0_RVT U2527 ( .A1(n2320), .A2(n1774), .Y(n580) );
  NAND2X0_RVT U2528 ( .A1(n2320), .A2(n1487), .Y(n573) );
  OA22X1_RVT U2529 ( .A1(n574), .A2(n1695), .A3(n573), .A4(n1816), .Y(n597) );
  AO221X1_RVT U2530 ( .A1(N974), .A2(net32868), .A3(N1031), .A4(net32878), 
        .A5(n1856), .Y(N1089) );
  OA22X1_RVT U2531 ( .A1(n577), .A2(n1695), .A3(n574), .A4(n1816), .Y(n589) );
  AO221X1_RVT U2532 ( .A1(N975), .A2(net32868), .A3(N1032), .A4(net32878), 
        .A5(n1015), .Y(N1090) );
  AO221X1_RVT U2533 ( .A1(N976), .A2(net32868), .A3(N1033), .A4(net32878), 
        .A5(n1015), .Y(N1091) );
  AO221X1_RVT U2534 ( .A1(N977), .A2(net32868), .A3(N1034), .A4(net32878), 
        .A5(n1015), .Y(N1092) );
  AO221X1_RVT U2535 ( .A1(N978), .A2(net32868), .A3(N1035), .A4(net32878), 
        .A5(n1015), .Y(N1093) );
  AO221X1_RVT U2536 ( .A1(N979), .A2(net32868), .A3(N1036), .A4(net32880), 
        .A5(n1015), .Y(N1094) );
  AO221X1_RVT U2537 ( .A1(N980), .A2(net32868), .A3(N1037), .A4(net32880), 
        .A5(n1015), .Y(N1095) );
  AO22X1_RVT U2538 ( .A1(N155), .A2(net32926), .A3(N464), .A4(net32958), .Y(
        n2107) );
  AO22X1_RVT U2539 ( .A1(N999), .A2(net32880), .A3(N942), .A4(net32866), .Y(
        n2104) );
  AO221X1_RVT U2540 ( .A1(N239), .A2(net32932), .A3(N213), .A4(net32938), .A5(
        n2104), .Y(n2105) );
  NAND3X0_RVT U2541 ( .A1(n1768), .A2(n1485), .A3(n1494), .Y(n2288) );
  NAND3X0_RVT U2542 ( .A1(n1768), .A2(n1494), .A3(n2288), .Y(n2294) );
  OA22X1_RVT U2543 ( .A1(n1825), .A2(n1695), .A3(n1815), .A4(n1816), .Y(n516)
         );
  AO221X1_RVT U2544 ( .A1(N981), .A2(net32868), .A3(N1038), .A4(net32880), 
        .A5(n1856), .Y(N1096) );
  AO22X1_RVT U2545 ( .A1(N154), .A2(net32926), .A3(N463), .A4(net32958), .Y(
        n2112) );
  AO222X1_RVT U2546 ( .A1(N438), .A2(net32946), .A3(N354), .A4(net32952), .A5(
        N412), .A6(net27438), .Y(n2111) );
  AO22X1_RVT U2547 ( .A1(N998), .A2(net32880), .A3(N941), .A4(net32866), .Y(
        n2109) );
  AO221X1_RVT U2548 ( .A1(N238), .A2(net32932), .A3(N212), .A4(net32938), .A5(
        n2109), .Y(n2110) );
  NAND2X0_RVT U2549 ( .A1(tmp_m0[4]), .A2(n2315), .Y(n426) );
  NAND2X0_RVT U2550 ( .A1(n2322), .A2(n2113), .Y(n461) );
  OA22X1_RVT U2551 ( .A1(n461), .A2(n1695), .A3(n1825), .A4(n1816), .Y(n502)
         );
  AO221X1_RVT U2552 ( .A1(N982), .A2(net32868), .A3(N1039), .A4(net32880), 
        .A5(n1856), .Y(N1097) );
  NAND2X0_RVT U2553 ( .A1(n2322), .A2(n2114), .Y(n464) );
  OA22X1_RVT U2554 ( .A1(n464), .A2(n1695), .A3(n461), .A4(n1816), .Y(n487) );
  AO221X1_RVT U2555 ( .A1(N983), .A2(net32870), .A3(N1040), .A4(net32880), 
        .A5(n1856), .Y(N1098) );
  AO22X1_RVT U2556 ( .A1(N152), .A2(net32926), .A3(N461), .A4(net32958), .Y(
        n2118) );
  AO222X1_RVT U2557 ( .A1(N436), .A2(net32946), .A3(N352), .A4(net32952), .A5(
        N410), .A6(net32962), .Y(n2117) );
  AO22X1_RVT U2558 ( .A1(N996), .A2(net32880), .A3(N939), .A4(net32866), .Y(
        n2115) );
  AO22X1_RVT U2559 ( .A1(N151), .A2(net32924), .A3(N460), .A4(net32958), .Y(
        n2122) );
  AO222X1_RVT U2560 ( .A1(N435), .A2(net32946), .A3(N351), .A4(net32952), .A5(
        N409), .A6(net27438), .Y(n2121) );
  AO22X1_RVT U2561 ( .A1(N995), .A2(net32882), .A3(N938), .A4(net32866), .Y(
        n2119) );
  AO221X1_RVT U2562 ( .A1(N235), .A2(net32930), .A3(N209), .A4(net32938), .A5(
        n2119), .Y(n2120) );
  NAND2X0_RVT U2563 ( .A1(n1462), .A2(n1778), .Y(n2123) );
  OA22X1_RVT U2564 ( .A1(n463), .A2(n1695), .A3(n464), .A4(n1816), .Y(n462) );
  MUX21X1_RVT U2565 ( .A1(b_m[22]), .A2(n1251), .S0(n1941), .Y(n1381) );
  MUX21X1_RVT U2566 ( .A1(n1938), .A2(n1250), .S0(n1942), .Y(n1379) );
  MUX21X1_RVT U2567 ( .A1(b_m[20]), .A2(n1249), .S0(n1941), .Y(n1377) );
  MUX21X1_RVT U2568 ( .A1(b_m[19]), .A2(n1248), .S0(n1942), .Y(n1375) );
  MUX21X1_RVT U2569 ( .A1(b_m[18]), .A2(n1247), .S0(n1940), .Y(n1373) );
  MUX21X1_RVT U2570 ( .A1(n1936), .A2(n1246), .S0(n1943), .Y(n1371) );
  MUX21X1_RVT U2571 ( .A1(n1934), .A2(n1245), .S0(n1941), .Y(n1369) );
  MUX21X1_RVT U2572 ( .A1(b_m[15]), .A2(n1244), .S0(n1940), .Y(n1367) );
  MUX21X1_RVT U2573 ( .A1(b_m[14]), .A2(n1243), .S0(n1941), .Y(n1365) );
  MUX21X1_RVT U2574 ( .A1(n1411), .A2(n1242), .S0(rst), .Y(n1363) );
  MUX21X1_RVT U2575 ( .A1(b_m[12]), .A2(n1241), .S0(n1940), .Y(n1361) );
  MUX21X1_RVT U2576 ( .A1(b_m[11]), .A2(n1240), .S0(n1943), .Y(n1359) );
  MUX21X1_RVT U2577 ( .A1(b_m[10]), .A2(n1239), .S0(n1942), .Y(n1357) );
  MUX21X1_RVT U2578 ( .A1(b_m[9]), .A2(n1238), .S0(n1943), .Y(n1355) );
  MUX21X1_RVT U2579 ( .A1(n1932), .A2(n1237), .S0(n1942), .Y(n1353) );
  MUX21X1_RVT U2580 ( .A1(b_m[7]), .A2(n1236), .S0(n1943), .Y(n1351) );
  MUX21X1_RVT U2581 ( .A1(b_m[6]), .A2(n1235), .S0(n1940), .Y(n1349) );
  MUX21X1_RVT U2582 ( .A1(n1931), .A2(n1234), .S0(n1944), .Y(n1347) );
  MUX21X1_RVT U2583 ( .A1(b_m[4]), .A2(n1233), .S0(n1940), .Y(n1345) );
  MUX21X1_RVT U2584 ( .A1(b_m[3]), .A2(n1232), .S0(n1944), .Y(n1343) );
  MUX21X1_RVT U2585 ( .A1(n1930), .A2(n1231), .S0(n1942), .Y(n1341) );
  MUX21X1_RVT U2586 ( .A1(b_m[1]), .A2(n1230), .S0(n1944), .Y(n1339) );
  MUX21X1_RVT U2587 ( .A1(n1928), .A2(n1229), .S0(n1940), .Y(n1337) );
  MUX21X1_RVT U2588 ( .A1(n1464), .A2(n1226), .S0(n1944), .Y(n1333) );
  MUX21X1_RVT U2589 ( .A1(n1505), .A2(n1225), .S0(n1942), .Y(n1331) );
  MUX21X1_RVT U2590 ( .A1(a_m[20]), .A2(n1224), .S0(n1945), .Y(n1329) );
  MUX21X1_RVT U2591 ( .A1(n1465), .A2(n1223), .S0(rst), .Y(n1327) );
  MUX21X1_RVT U2592 ( .A1(n1506), .A2(n1222), .S0(n1945), .Y(n1325) );
  MUX21X1_RVT U2593 ( .A1(n1472), .A2(n1221), .S0(n1941), .Y(n1323) );
  MUX21X1_RVT U2594 ( .A1(n1488), .A2(n1220), .S0(n1945), .Y(n1321) );
  MUX21X1_RVT U2595 ( .A1(n1460), .A2(n1219), .S0(rst), .Y(n1319) );
  MUX21X1_RVT U2596 ( .A1(n1507), .A2(n1218), .S0(n1945), .Y(n1317) );
  MUX21X1_RVT U2597 ( .A1(n1489), .A2(n1217), .S0(n1943), .Y(n1315) );
  MUX21X1_RVT U2598 ( .A1(n1508), .A2(n1216), .S0(n1945), .Y(n1313) );
  MUX21X1_RVT U2599 ( .A1(a_m[11]), .A2(n1215), .S0(n1941), .Y(n1311) );
  MUX21X1_RVT U2600 ( .A1(n1481), .A2(n1214), .S0(n1945), .Y(n1309) );
  MUX21X1_RVT U2601 ( .A1(a_m[9]), .A2(n1213), .S0(n1943), .Y(n1307) );
  MUX21X1_RVT U2602 ( .A1(n1480), .A2(n1212), .S0(rst), .Y(n1305) );
  MUX21X1_RVT U2603 ( .A1(n1466), .A2(n1211), .S0(n1943), .Y(n1303) );
  MUX21X1_RVT U2604 ( .A1(n1509), .A2(n1210), .S0(n1946), .Y(n1301) );
  MUX21X1_RVT U2605 ( .A1(n1482), .A2(n1209), .S0(n1942), .Y(n1299) );
  MUX21X1_RVT U2606 ( .A1(n1510), .A2(n1208), .S0(n1946), .Y(n1297) );
  MUX21X1_RVT U2607 ( .A1(n1483), .A2(n1207), .S0(n1944), .Y(n1295) );
  MUX21X1_RVT U2608 ( .A1(n1490), .A2(n1206), .S0(n1946), .Y(n1293) );
  MUX21X1_RVT U2609 ( .A1(n1511), .A2(n1205), .S0(n1944), .Y(n1291) );
  MUX21X1_RVT U2610 ( .A1(a_m[0]), .A2(n1204), .S0(n1946), .Y(n1289) );
  MUX21X1_RVT U2611 ( .A1(n1871), .A2(n1471), .S0(N1129), .Y(n2125) );
  AO21X1_RVT U2612 ( .A1(N1886), .A2(tmp_m0[24]), .A3(n2125), .Y(n1007) );
  NAND4X0_RVT U2613 ( .A1(n1593), .A2(n2289), .A3(n1478), .A4(n2287), .Y(n1002) );
  AO222X1_RVT U2614 ( .A1(N1670), .A2(n1871), .A3(n1910), .A4(n1471), .A5(
        N1887), .A6(tmp_m0[24]), .Y(n982) );
  OA22X1_RVT U2615 ( .A1(n1870), .A2(n1816), .A3(n1486), .A4(n1843), .Y(n625)
         );
  OA22X1_RVT U2616 ( .A1(n1881), .A2(n1695), .A3(n1504), .A4(n1885), .Y(n627)
         );
  OA222X1_RVT U2617 ( .A1(n1881), .A2(n1816), .A3(n1690), .A4(n1886), .A5(
        n1475), .A6(n1868), .Y(n621) );
  OA222X1_RVT U2618 ( .A1(n1702), .A2(n1695), .A3(n1504), .A4(n1860), .A5(
        n2316), .A6(n1892), .Y(n622) );
  OA22X1_RVT U2619 ( .A1(n2316), .A2(n1869), .A3(n1623), .A4(n1843), .Y(n612)
         );
  OA222X1_RVT U2620 ( .A1(n1818), .A2(n1695), .A3(n1690), .A4(n1860), .A5(
        n1702), .A6(n1816), .Y(n615) );
  OA22X1_RVT U2621 ( .A1(n1504), .A2(n1869), .A3(n1787), .A4(n1843), .Y(n606)
         );
  OA222X1_RVT U2622 ( .A1(n580), .A2(n1695), .A3(n1475), .A4(n1702), .A5(n1818), .A6(n1816), .Y(n609) );
  OA222X1_RVT U2623 ( .A1(n1690), .A2(n1869), .A3(n1789), .A4(n1844), .A5(
        n1787), .A6(n1873), .Y(n600) );
  OA222X1_RVT U2624 ( .A1(n573), .A2(n1695), .A3(n1475), .A4(n1818), .A5(n580), 
        .A6(n1816), .Y(n603) );
  OA222X1_RVT U2625 ( .A1(n1545), .A2(n1869), .A3(n1496), .A4(n1844), .A5(
        n1789), .A6(n1873), .Y(n593) );
  OA222X1_RVT U2626 ( .A1(n1486), .A2(n1869), .A3(n1520), .A4(n1844), .A5(
        n1496), .A6(n1873), .Y(n585) );
  OA222X1_RVT U2627 ( .A1(n1470), .A2(n1869), .A3(n1476), .A4(n1844), .A5(
        n1520), .A6(n1873), .Y(n569) );
  OA22X1_RVT U2628 ( .A1(n2316), .A2(n1821), .A3(n1486), .A4(n1842), .Y(n563)
         );
  OA22X1_RVT U2629 ( .A1(n1802), .A2(n1695), .A3(n1475), .A4(n408), .Y(n565)
         );
  OA22X1_RVT U2630 ( .A1(n1824), .A2(n1816), .A3(n1545), .A4(n402), .Y(n566)
         );
  OA22X1_RVT U2631 ( .A1(n1623), .A2(n1869), .A3(n1461), .A4(n1843), .Y(n558)
         );
  OA22X1_RVT U2632 ( .A1(n1787), .A2(n1869), .A3(n1612), .A4(n1843), .Y(n547)
         );
  NAND2X0_RVT U2633 ( .A1(n1544), .A2(tmp_m0[29]), .Y(n2127) );
  OA222X1_RVT U2634 ( .A1(n1470), .A2(n1842), .A3(n1802), .A4(n1816), .A5(
        n2316), .A6(n408), .Y(n2126) );
  AND4X1_RVT U2635 ( .A1(n553), .A2(n555), .A3(n2127), .A4(n2126), .Y(n2128)
         );
  OA222X1_RVT U2636 ( .A1(n648), .A2(n2128), .A3(n1496), .A4(n1860), .A5(n1786), .A6(n1695), .Y(n550) );
  OA22X1_RVT U2637 ( .A1(n1789), .A2(n1869), .A3(n1611), .A4(n1843), .Y(n536)
         );
  OA22X1_RVT U2638 ( .A1(n1690), .A2(n1821), .A3(n1623), .A4(n1842), .Y(n2129)
         );
  OA222X1_RVT U2639 ( .A1(n648), .A2(n2130), .A3(n1811), .A4(n1816), .A5(n1805), .A6(n1695), .Y(n539) );
  OA22X1_RVT U2640 ( .A1(n1545), .A2(n1821), .A3(n1787), .A4(n1842), .Y(n530)
         );
  OA222X1_RVT U2641 ( .A1(n1496), .A2(n1869), .A3(n1615), .A4(n1844), .A5(
        n1611), .A6(n1873), .Y(n525) );
  OA222X1_RVT U2642 ( .A1(n1815), .A2(n1695), .A3(n1475), .A4(n1810), .A5(
        n1805), .A6(n1816), .Y(n528) );
  OA22X1_RVT U2643 ( .A1(n1486), .A2(n1821), .A3(n1789), .A4(n1842), .Y(n519)
         );
  OA222X1_RVT U2644 ( .A1(n1520), .A2(n1868), .A3(n1795), .A4(n1559), .A5(
        n1615), .A6(n1873), .Y(n511) );
  OA22X1_RVT U2645 ( .A1(n1470), .A2(n1821), .A3(n1496), .A4(n1792), .Y(n504)
         );
  OA22X1_RVT U2646 ( .A1(n1623), .A2(n1821), .A3(n1520), .A4(n1842), .Y(n490)
         );
  OA222X1_RVT U2647 ( .A1(n1461), .A2(n1868), .A3(n1606), .A4(n1559), .A5(
        n1625), .A6(n1873), .Y(n482) );
  OA22X1_RVT U2648 ( .A1(n1787), .A2(n1821), .A3(n1476), .A4(n1842), .Y(n470)
         );
  OA22X1_RVT U2649 ( .A1(n1561), .A2(n1844), .A3(n1612), .A4(n1868), .Y(n2131)
         );
  OA221X1_RVT U2650 ( .A1(n1606), .A2(n1874), .A3(n1625), .A4(n1876), .A5(
        n2131), .Y(n456) );
  OA22X1_RVT U2651 ( .A1(n1690), .A2(n2293), .A3(n1486), .A4(n2301), .Y(n418)
         );
  OA22X1_RVT U2652 ( .A1(n432), .A2(n1695), .A3(n1504), .A4(n2294), .Y(n419)
         );
  OA22X1_RVT U2653 ( .A1(n2290), .A2(n1816), .A3(n1545), .A4(n2295), .Y(n421)
         );
  OA22X1_RVT U2654 ( .A1(n1789), .A2(n1821), .A3(n1461), .A4(n1842), .Y(n398)
         );
  AO22X1_RVT U2655 ( .A1(N459), .A2(net32958), .A3(N408), .A4(net27438), .Y(
        n2136) );
  AO22X1_RVT U2656 ( .A1(N434), .A2(net32946), .A3(N350), .A4(net32952), .Y(
        n2135) );
  AO22X1_RVT U2657 ( .A1(N937), .A2(net32870), .A3(N208), .A4(net27434), .Y(
        n2133) );
  AO221X1_RVT U2658 ( .A1(N150), .A2(net32924), .A3(N234), .A4(net32930), .A5(
        n2133), .Y(n2134) );
  OR3X1_RVT U2659 ( .A1(n2136), .A2(n2135), .A3(n2134), .Y(n2137) );
  AO21X1_RVT U2660 ( .A1(N994), .A2(net32882), .A3(n2137), .Y(N1052) );
  AO22X1_RVT U2661 ( .A1(tmp_m0[1]), .A2(n619), .A3(tmp_m0[0]), .A4(n620), .Y(
        N2065) );
  AO222X1_RVT U2662 ( .A1(tmp_m0[1]), .A2(n620), .A3(tmp_m0[2]), .A4(n619), 
        .A5(tmp_m0[0]), .A6(n617), .Y(N2066) );
  AO22X1_RVT U2663 ( .A1(tmp_m0[1]), .A2(n617), .A3(tmp_m0[2]), .A4(n620), .Y(
        n2138) );
  AO221X1_RVT U2664 ( .A1(n2153), .A2(tmp_m0[0]), .A3(tmp_m0[3]), .A4(n619), 
        .A5(n2138), .Y(N2067) );
  NAND2X0_RVT U2665 ( .A1(n619), .A2(tmp_m0[4]), .Y(n2141) );
  AOI22X1_RVT U2666 ( .A1(tmp_m0[2]), .A2(n617), .A3(n620), .A4(tmp_m0[3]), 
        .Y(n2140) );
  NAND4X0_RVT U2667 ( .A1(n2143), .A2(n2142), .A3(n2141), .A4(n2140), .Y(N2068) );
  AO222X1_RVT U2668 ( .A1(tmp_m0[2]), .A2(n1890), .A3(tmp_m0[1]), .A4(n1863), 
        .A5(tmp_m0[0]), .A6(n1899), .Y(n2145) );
  AO22X1_RVT U2669 ( .A1(tmp_m0[3]), .A2(n617), .A3(tmp_m0[4]), .A4(n620), .Y(
        n2144) );
  AO221X1_RVT U2670 ( .A1(n2145), .A2(n1852), .A3(tmp_m0[5]), .A4(n619), .A5(
        n2144), .Y(N2069) );
  AO22X1_RVT U2671 ( .A1(tmp_m0[1]), .A2(n1900), .A3(tmp_m0[3]), .A4(n1890), 
        .Y(n2146) );
  AO221X1_RVT U2672 ( .A1(tmp_m0[2]), .A2(n1863), .A3(tmp_m0[0]), .A4(n1871), 
        .A5(n2146), .Y(n2148) );
  AO22X1_RVT U2673 ( .A1(tmp_m0[4]), .A2(n617), .A3(tmp_m0[5]), .A4(n620), .Y(
        n2147) );
  NAND4X0_RVT U2674 ( .A1(n643), .A2(n644), .A3(n1861), .A4(n2149), .Y(n2151)
         );
  AO22X1_RVT U2675 ( .A1(n1866), .A2(tmp_m0[24]), .A3(n1846), .A4(tmp_m0[22]), 
        .Y(n2150) );
  AO221X1_RVT U2676 ( .A1(n2151), .A2(n1852), .A3(tmp_m0[23]), .A4(n1858), 
        .A5(n2150), .Y(N2088) );
  AO22X1_RVT U2677 ( .A1(tmp_m0[25]), .A2(n619), .A3(tmp_m0[24]), .A4(n1859), 
        .Y(N2089) );
  AO222X1_RVT U2678 ( .A1(tmp_m0[25]), .A2(n620), .A3(tmp_m0[26]), .A4(n619), 
        .A5(n1845), .A6(tmp_m0[24]), .Y(N2090) );
  AO222X1_RVT U2679 ( .A1(tmp_m0[26]), .A2(n620), .A3(n619), .A4(tmp_m0[27]), 
        .A5(tmp_m0[25]), .A6(n617), .Y(N2091) );
  AO22X1_RVT U2680 ( .A1(tmp_m0[26]), .A2(n617), .A3(n620), .A4(tmp_m0[27]), 
        .Y(n2152) );
  AO221X1_RVT U2681 ( .A1(tmp_m0[25]), .A2(n2153), .A3(n619), .A4(tmp_m0[28]), 
        .A5(n2152), .Y(N2092) );
  OA22X1_RVT U2682 ( .A1(n1861), .A2(n2291), .A3(n1873), .A4(n1494), .Y(n2157)
         );
  OA22X1_RVT U2683 ( .A1(n1869), .A2(n1462), .A3(n1879), .A4(n1533), .Y(n2156)
         );
  OA22X1_RVT U2684 ( .A1(n1877), .A2(n1485), .A3(n1885), .A4(n1497), .Y(n2155)
         );
  OA22X1_RVT U2685 ( .A1(n1893), .A2(n2287), .A3(n1813), .A4(n1843), .Y(n2154)
         );
  NAND4X0_RVT U2686 ( .A1(n2157), .A2(n2156), .A3(n2155), .A4(n2154), .Y(n2159) );
  AO22X1_RVT U2687 ( .A1(n1866), .A2(tmp_m0[7]), .A3(n1846), .A4(tmp_m0[5]), 
        .Y(n2158) );
  AO221X1_RVT U2688 ( .A1(n2159), .A2(n1852), .A3(tmp_m0[6]), .A4(n1858), .A5(
        n2158), .Y(N2071) );
  OA222X1_RVT U2689 ( .A1(n1874), .A2(n1813), .A3(n1702), .A4(n1533), .A5(
        n1861), .A6(n1497), .Y(n2163) );
  OA22X1_RVT U2690 ( .A1(n1870), .A2(n1778), .A3(n1879), .A4(n2289), .Y(n2162)
         );
  OA22X1_RVT U2691 ( .A1(n1877), .A2(n1494), .A3(n1885), .A4(n1485), .Y(n2161)
         );
  OA22X1_RVT U2692 ( .A1(n1893), .A2(n2291), .A3(n2301), .A4(n1559), .Y(n2160)
         );
  NAND4X0_RVT U2693 ( .A1(n2163), .A2(n2162), .A3(n2161), .A4(n2160), .Y(n2165) );
  AO22X1_RVT U2694 ( .A1(n1866), .A2(tmp_m0[8]), .A3(n1846), .A4(tmp_m0[6]), 
        .Y(n2164) );
  AO221X1_RVT U2695 ( .A1(n2165), .A2(n1852), .A3(tmp_m0[7]), .A4(n1858), .A5(
        n2164), .Y(N2072) );
  OA222X1_RVT U2696 ( .A1(n1874), .A2(n2301), .A3(n1702), .A4(n2289), .A5(
        n1861), .A6(n1485), .Y(n2169) );
  OA22X1_RVT U2697 ( .A1(n1869), .A2(n2291), .A3(n1879), .A4(n2287), .Y(n2168)
         );
  OA222X1_RVT U2698 ( .A1(n1818), .A2(n1533), .A3(n1876), .A4(n1813), .A5(
        n1885), .A6(n1494), .Y(n2167) );
  OA22X1_RVT U2699 ( .A1(n1893), .A2(n1497), .A3(n1803), .A4(n1559), .Y(n2166)
         );
  NAND4X0_RVT U2700 ( .A1(n2169), .A2(n2168), .A3(n2167), .A4(n2166), .Y(n2171) );
  AO22X1_RVT U2701 ( .A1(n1866), .A2(tmp_m0[9]), .A3(n1846), .A4(tmp_m0[7]), 
        .Y(n2170) );
  AO221X1_RVT U2702 ( .A1(n2171), .A2(n1852), .A3(tmp_m0[8]), .A4(n1858), .A5(
        n2170), .Y(N2073) );
  OA222X1_RVT U2703 ( .A1(n1874), .A2(n1803), .A3(n1702), .A4(n2287), .A5(
        n1861), .A6(n1494), .Y(n2175) );
  OA222X1_RVT U2704 ( .A1(n1876), .A2(n2301), .A3(n1868), .A4(n1497), .A5(
        n1879), .A6(n2291), .Y(n2174) );
  OA222X1_RVT U2705 ( .A1(n580), .A2(n1533), .A3(n1885), .A4(n1813), .A5(n1818), .A6(n2289), .Y(n2173) );
  OA22X1_RVT U2706 ( .A1(n1893), .A2(n1485), .A3(n1469), .A4(n1559), .Y(n2172)
         );
  NAND4X0_RVT U2707 ( .A1(n2175), .A2(n2174), .A3(n2173), .A4(n2172), .Y(n2177) );
  AO22X1_RVT U2708 ( .A1(n1866), .A2(tmp_m0[10]), .A3(n1846), .A4(tmp_m0[8]), 
        .Y(n2176) );
  AO221X1_RVT U2709 ( .A1(n2177), .A2(n1852), .A3(tmp_m0[9]), .A4(n1858), .A5(
        n2176), .Y(N2074) );
  OA222X1_RVT U2710 ( .A1(n1801), .A2(n1559), .A3(n580), .A4(n2289), .A5(n1892), .A6(n1494), .Y(n2178) );
  AO22X1_RVT U2711 ( .A1(n1866), .A2(tmp_m0[11]), .A3(n1846), .A4(tmp_m0[9]), 
        .Y(n2179) );
  OA22X1_RVT U2712 ( .A1(n1873), .A2(n1801), .A3(n1868), .A4(n1494), .Y(n2181)
         );
  OA222X1_RVT U2713 ( .A1(n1473), .A2(n1559), .A3(n580), .A4(n1778), .A5(n1892), .A6(n1813), .Y(n2182) );
  AO22X1_RVT U2714 ( .A1(n1866), .A2(tmp_m0[12]), .A3(n1846), .A4(tmp_m0[10]), 
        .Y(n2183) );
  OA22X1_RVT U2715 ( .A1(n1873), .A2(n1473), .A3(n1868), .A4(n1813), .Y(n2185)
         );
  OA221X1_RVT U2716 ( .A1(n1860), .A2(n1803), .A3(n1702), .A4(n1485), .A5(
        n2185), .Y(n2190) );
  OA222X1_RVT U2717 ( .A1(n1886), .A2(n1469), .A3(n1880), .A4(n1494), .A5(
        n1875), .A6(n1801), .Y(n2189) );
  OA22X1_RVT U2718 ( .A1(n574), .A2(n1462), .A3(n573), .A4(n2287), .Y(n2186)
         );
  OA221X1_RVT U2719 ( .A1(n577), .A2(n1533), .A3(n1818), .A4(n1497), .A5(n2186), .Y(n2188) );
  OA222X1_RVT U2720 ( .A1(n1613), .A2(n1559), .A3(n580), .A4(n2291), .A5(n1892), .A6(n2301), .Y(n2187) );
  AO22X1_RVT U2721 ( .A1(n1866), .A2(tmp_m0[13]), .A3(n1846), .A4(tmp_m0[11]), 
        .Y(n2191) );
  OA22X1_RVT U2722 ( .A1(n1873), .A2(n1613), .A3(n1868), .A4(n2301), .Y(n2193)
         );
  OA22X1_RVT U2723 ( .A1(n1887), .A2(n1801), .A3(n1818), .A4(n1485), .Y(n2194)
         );
  OA22X1_RVT U2724 ( .A1(n574), .A2(n2287), .A3(n573), .A4(n2291), .Y(n2195)
         );
  AO22X1_RVT U2725 ( .A1(n1866), .A2(tmp_m0[14]), .A3(n1847), .A4(tmp_m0[12]), 
        .Y(n2197) );
  AO221X1_RVT U2726 ( .A1(n2198), .A2(n1560), .A3(tmp_m0[13]), .A4(n1858), 
        .A5(n2197), .Y(N2078) );
  OA22X1_RVT U2727 ( .A1(n2291), .A2(n1821), .A3(n1822), .A4(n1497), .Y(n2202)
         );
  OA22X1_RVT U2728 ( .A1(n1819), .A2(n1485), .A3(n1802), .A4(n1533), .Y(n2201)
         );
  OA22X1_RVT U2729 ( .A1(n408), .A2(n2287), .A3(n402), .A4(n1494), .Y(n2200)
         );
  OA22X1_RVT U2730 ( .A1(n1824), .A2(n2289), .A3(n1813), .A4(n1842), .Y(n2199)
         );
  AND4X1_RVT U2731 ( .A1(n2202), .A2(n2201), .A3(n2200), .A4(n2199), .Y(n2203)
         );
  OA222X1_RVT U2732 ( .A1(n1874), .A2(n1790), .A3(n648), .A4(n2203), .A5(n1861), .A6(n1801), .Y(n2207) );
  OA22X1_RVT U2733 ( .A1(n1870), .A2(n1803), .A3(n1879), .A4(n2301), .Y(n2206)
         );
  OA22X1_RVT U2734 ( .A1(n1877), .A2(n1613), .A3(n1885), .A4(n1473), .Y(n2205)
         );
  OA22X1_RVT U2735 ( .A1(n1893), .A2(n1469), .A3(n1791), .A4(n1843), .Y(n2204)
         );
  NAND4X0_RVT U2736 ( .A1(n2207), .A2(n2206), .A3(n2205), .A4(n2204), .Y(n2209) );
  AO22X1_RVT U2737 ( .A1(n1866), .A2(tmp_m0[15]), .A3(n1846), .A4(tmp_m0[13]), 
        .Y(n2208) );
  AO221X1_RVT U2738 ( .A1(n2209), .A2(n1852), .A3(tmp_m0[14]), .A4(n1858), 
        .A5(n2208), .Y(N2079) );
  OA22X1_RVT U2739 ( .A1(n1497), .A2(n1821), .A3(n1822), .A4(n1485), .Y(n2213)
         );
  OA22X1_RVT U2740 ( .A1(n1819), .A2(n1494), .A3(n1802), .A4(n1462), .Y(n2212)
         );
  OA22X1_RVT U2741 ( .A1(n408), .A2(n2291), .A3(n402), .A4(n1813), .Y(n2211)
         );
  OA22X1_RVT U2742 ( .A1(n1824), .A2(n2287), .A3(n2301), .A4(n1842), .Y(n2210)
         );
  AND4X1_RVT U2743 ( .A1(n2213), .A2(n2212), .A3(n2211), .A4(n2210), .Y(n2214)
         );
  OA222X1_RVT U2744 ( .A1(n1860), .A2(n1473), .A3(n648), .A4(n2214), .A5(n1786), .A6(n1533), .Y(n2218) );
  OA22X1_RVT U2745 ( .A1(n1874), .A2(n1791), .A3(n1868), .A4(n1469), .Y(n2217)
         );
  OA222X1_RVT U2746 ( .A1(n1886), .A2(n1613), .A3(n1880), .A4(n1803), .A5(
        n1875), .A6(n1790), .Y(n2216) );
  OA22X1_RVT U2747 ( .A1(n1893), .A2(n1801), .A3(n1842), .A4(n1843), .Y(n2215)
         );
  AO22X1_RVT U2748 ( .A1(n1866), .A2(tmp_m0[16]), .A3(n1846), .A4(tmp_m0[14]), 
        .Y(n2219) );
  AO221X1_RVT U2749 ( .A1(n2220), .A2(n1852), .A3(tmp_m0[15]), .A4(n1859), 
        .A5(n2219), .Y(N2080) );
  OA22X1_RVT U2750 ( .A1(n1485), .A2(n1821), .A3(n1822), .A4(n1494), .Y(n2224)
         );
  OA22X1_RVT U2751 ( .A1(n1819), .A2(n1813), .A3(n1802), .A4(n2287), .Y(n2223)
         );
  OA22X1_RVT U2752 ( .A1(n408), .A2(n1497), .A3(n402), .A4(n2301), .Y(n2222)
         );
  OA22X1_RVT U2753 ( .A1(n1824), .A2(n2291), .A3(n1803), .A4(n1842), .Y(n2221)
         );
  AND4X1_RVT U2754 ( .A1(n2224), .A2(n2223), .A3(n2222), .A4(n2221), .Y(n2225)
         );
  OA222X1_RVT U2755 ( .A1(n1806), .A2(n1533), .A3(n648), .A4(n2225), .A5(n1786), .A6(n2289), .Y(n2229) );
  OA222X1_RVT U2756 ( .A1(n1869), .A2(n1801), .A3(n1860), .A4(n1613), .A5(
        n1873), .A6(n1842), .Y(n2228) );
  OA222X1_RVT U2757 ( .A1(n1886), .A2(n1790), .A3(n1880), .A4(n1469), .A5(
        n1875), .A6(n1791), .Y(n2227) );
  OA22X1_RVT U2758 ( .A1(n1893), .A2(n1473), .A3(n1468), .A4(n1843), .Y(n2226)
         );
  AO22X1_RVT U2759 ( .A1(n1866), .A2(tmp_m0[17]), .A3(n1846), .A4(tmp_m0[15]), 
        .Y(n2230) );
  AO221X1_RVT U2760 ( .A1(n2231), .A2(n1852), .A3(tmp_m0[16]), .A4(n1859), 
        .A5(n2230), .Y(N2081) );
  OA22X1_RVT U2761 ( .A1(n1494), .A2(n1821), .A3(n1822), .A4(n1813), .Y(n2235)
         );
  OA22X1_RVT U2762 ( .A1(n1819), .A2(n2301), .A3(n1802), .A4(n2291), .Y(n2234)
         );
  OA22X1_RVT U2763 ( .A1(n408), .A2(n1485), .A3(n402), .A4(n1803), .Y(n2233)
         );
  OA22X1_RVT U2764 ( .A1(n1824), .A2(n1497), .A3(n1469), .A4(n1842), .Y(n2232)
         );
  AND4X1_RVT U2765 ( .A1(n2235), .A2(n2234), .A3(n2233), .A4(n2232), .Y(n2236)
         );
  OA222X1_RVT U2766 ( .A1(n1484), .A2(n1559), .A3(n1885), .A4(n1791), .A5(
        n1892), .A6(n1613), .Y(n2237) );
  AO22X1_RVT U2767 ( .A1(n1866), .A2(tmp_m0[18]), .A3(n1846), .A4(tmp_m0[16]), 
        .Y(n2238) );
  OA22X1_RVT U2768 ( .A1(n1813), .A2(n1821), .A3(n1822), .A4(n2301), .Y(n2243)
         );
  OA22X1_RVT U2769 ( .A1(n1819), .A2(n1803), .A3(n1802), .A4(n1497), .Y(n2242)
         );
  OA22X1_RVT U2770 ( .A1(n408), .A2(n1494), .A3(n402), .A4(n1469), .Y(n2241)
         );
  OA22X1_RVT U2771 ( .A1(n1824), .A2(n1485), .A3(n1801), .A4(n1842), .Y(n2240)
         );
  AND4X1_RVT U2772 ( .A1(n2243), .A2(n2242), .A3(n2241), .A4(n2240), .Y(n2245)
         );
  OA22X1_RVT U2773 ( .A1(n1806), .A2(n2287), .A3(n1815), .A4(n2289), .Y(n2244)
         );
  OA222X1_RVT U2774 ( .A1(n1492), .A2(n1559), .A3(n1825), .A4(n1533), .A5(
        n1892), .A6(n1790), .Y(n2246) );
  AO22X1_RVT U2775 ( .A1(n1866), .A2(tmp_m0[19]), .A3(n1846), .A4(tmp_m0[17]), 
        .Y(n2247) );
  OA22X1_RVT U2776 ( .A1(n2301), .A2(n1821), .A3(n1822), .A4(n1803), .Y(n2252)
         );
  OA22X1_RVT U2777 ( .A1(n1819), .A2(n1469), .A3(n1802), .A4(n1485), .Y(n2251)
         );
  OA22X1_RVT U2778 ( .A1(n408), .A2(n1813), .A3(n402), .A4(n1801), .Y(n2250)
         );
  OA22X1_RVT U2779 ( .A1(n1824), .A2(n1494), .A3(n1473), .A4(n1842), .Y(n2249)
         );
  AND4X1_RVT U2780 ( .A1(n2252), .A2(n2251), .A3(n2250), .A4(n2249), .Y(n2254)
         );
  OA22X1_RVT U2781 ( .A1(n1806), .A2(n2291), .A3(n1815), .A4(n2287), .Y(n2253)
         );
  OA221X1_RVT U2782 ( .A1(n1692), .A2(n1497), .A3(n648), .A4(n2254), .A5(n2253), .Y(n2258) );
  OA222X1_RVT U2783 ( .A1(n1869), .A2(n1790), .A3(n1860), .A4(n1842), .A5(
        n1873), .A6(n1492), .Y(n2257) );
  OA22X1_RVT U2784 ( .A1(n1887), .A2(n1468), .A3(n461), .A4(n1533), .Y(n2255)
         );
  OA221X1_RVT U2785 ( .A1(n1877), .A2(n1484), .A3(n1880), .A4(n1613), .A5(
        n2255), .Y(n2256) );
  NAND4X0_RVT U2786 ( .A1(n2258), .A2(n2257), .A3(n2256), .A4(n1590), .Y(n2260) );
  AO22X1_RVT U2787 ( .A1(n1866), .A2(tmp_m0[20]), .A3(n1846), .A4(tmp_m0[18]), 
        .Y(n2259) );
  AO221X1_RVT U2788 ( .A1(n2260), .A2(n1851), .A3(tmp_m0[19]), .A4(n1859), 
        .A5(n2259), .Y(N2084) );
  OA22X1_RVT U2789 ( .A1(n1821), .A2(n1803), .A3(n1822), .A4(n1469), .Y(n2264)
         );
  OA22X1_RVT U2790 ( .A1(n1819), .A2(n1801), .A3(n1802), .A4(n1494), .Y(n2263)
         );
  OA22X1_RVT U2791 ( .A1(n408), .A2(n2301), .A3(n402), .A4(n1473), .Y(n2262)
         );
  OA22X1_RVT U2792 ( .A1(n1824), .A2(n1813), .A3(n1613), .A4(n1842), .Y(n2261)
         );
  AND4X1_RVT U2793 ( .A1(n2264), .A2(n2263), .A3(n2262), .A4(n2261), .Y(n2266)
         );
  OA22X1_RVT U2794 ( .A1(n1806), .A2(n1497), .A3(n1815), .A4(n2291), .Y(n2265)
         );
  OA22X1_RVT U2795 ( .A1(n1870), .A2(n1791), .A3(n1879), .A4(n1790), .Y(n2267)
         );
  OA22X1_RVT U2796 ( .A1(n464), .A2(n1533), .A3(n461), .A4(n2289), .Y(n2268)
         );
  OA222X1_RVT U2797 ( .A1(n1493), .A2(n1559), .A3(n1825), .A4(n1778), .A5(
        n1892), .A6(n1842), .Y(n2269) );
  AO22X1_RVT U2798 ( .A1(n1866), .A2(tmp_m0[21]), .A3(n1847), .A4(tmp_m0[19]), 
        .Y(n2270) );
  AO221X1_RVT U2799 ( .A1(n2271), .A2(n1851), .A3(tmp_m0[20]), .A4(n1859), 
        .A5(n2270), .Y(N2085) );
  OA22X1_RVT U2800 ( .A1(n1821), .A2(n1469), .A3(n1822), .A4(n1801), .Y(n2275)
         );
  OA22X1_RVT U2801 ( .A1(n1819), .A2(n1473), .A3(n1802), .A4(n1813), .Y(n2274)
         );
  OA22X1_RVT U2802 ( .A1(n408), .A2(n1803), .A3(n402), .A4(n1613), .Y(n2273)
         );
  OA22X1_RVT U2803 ( .A1(n1824), .A2(n2301), .A3(n1790), .A4(n1842), .Y(n2272)
         );
  AND4X1_RVT U2804 ( .A1(n2275), .A2(n2274), .A3(n2273), .A4(n2272), .Y(n2277)
         );
  OA22X1_RVT U2805 ( .A1(n1806), .A2(n1485), .A3(n1815), .A4(n1497), .Y(n2276)
         );
  OA221X1_RVT U2806 ( .A1(n1786), .A2(n1494), .A3(n648), .A4(n2277), .A5(n2276), .Y(n2284) );
  OA22X1_RVT U2807 ( .A1(n1870), .A2(n1842), .A3(n1879), .A4(n1791), .Y(n2278)
         );
  OA221X1_RVT U2808 ( .A1(n1874), .A2(n1493), .A3(n1861), .A4(n1484), .A5(
        n2278), .Y(n2283) );
  OA22X1_RVT U2809 ( .A1(n463), .A2(n1533), .A3(n464), .A4(n1462), .Y(n2279)
         );
  OA221X1_RVT U2810 ( .A1(n1887), .A2(n1492), .A3(n1875), .A4(n1518), .A5(
        n2279), .Y(n2282) );
  OA22X1_RVT U2811 ( .A1(n1893), .A2(n1468), .A3(n1474), .A4(n1843), .Y(n2280)
         );
  OA221X1_RVT U2812 ( .A1(n1825), .A2(n2291), .A3(n461), .A4(n1778), .A5(n2280), .Y(n2281) );
  AO22X1_RVT U2813 ( .A1(n1865), .A2(tmp_m0[22]), .A3(n1847), .A4(tmp_m0[20]), 
        .Y(n2285) );
  AO221X1_RVT U2814 ( .A1(n2286), .A2(n1851), .A3(tmp_m0[21]), .A4(n1859), 
        .A5(n2285), .Y(N2086) );
  OA21X1_RVT U2815 ( .A1(n2288), .A2(n1778), .A3(n426), .Y(n2292) );
  OA22X1_RVT U2816 ( .A1(n2292), .A2(n2291), .A3(n2290), .A4(n2289), .Y(n2299)
         );
  OA22X1_RVT U2817 ( .A1(n1497), .A2(n2294), .A3(n2293), .A4(n1485), .Y(n2298)
         );
  OA222X1_RVT U2818 ( .A1(n1813), .A2(n2301), .A3(n1494), .A4(n2295), .A5(n432), .A6(n1533), .Y(n2297) );
  NAND3X0_RVT U2819 ( .A1(n2299), .A2(n2298), .A3(n2297), .Y(n2308) );
  OA22X1_RVT U2820 ( .A1(n1821), .A2(n1801), .A3(n1822), .A4(n1473), .Y(n2306)
         );
  OA22X1_RVT U2821 ( .A1(n1819), .A2(n1613), .A3(n1802), .A4(n2301), .Y(n2305)
         );
  OA22X1_RVT U2822 ( .A1(n408), .A2(n1469), .A3(n402), .A4(n1790), .Y(n2304)
         );
  OA22X1_RVT U2823 ( .A1(n1824), .A2(n1803), .A3(n1791), .A4(n1842), .Y(n2303)
         );
  NAND4X0_RVT U2824 ( .A1(n2306), .A2(n2305), .A3(n2304), .A4(n2303), .Y(n2307) );
  AOI222X1_RVT U2825 ( .A1(tmp_m0[19]), .A2(n1863), .A3(n2308), .A4(n2322), 
        .A5(n2307), .A6(n2320), .Y(n2312) );
  OA22X1_RVT U2826 ( .A1(n1873), .A2(n1474), .A3(n1868), .A4(n1468), .Y(n2311)
         );
  OA222X1_RVT U2827 ( .A1(n1886), .A2(n1518), .A3(n1880), .A4(n1842), .A5(
        n1875), .A6(n1493), .Y(n2310) );
  OA22X1_RVT U2828 ( .A1(n1893), .A2(n1484), .A3(n1585), .A4(n1843), .Y(n2309)
         );
  NAND4X0_RVT U2829 ( .A1(n2312), .A2(n2311), .A3(n2310), .A4(n2309), .Y(n2314) );
  AO22X1_RVT U2830 ( .A1(n1865), .A2(tmp_m0[23]), .A3(n1847), .A4(tmp_m0[21]), 
        .Y(n2313) );
  AO221X1_RVT U2831 ( .A1(n2314), .A2(n1851), .A3(tmp_m0[22]), .A4(n1858), 
        .A5(n2313), .Y(N2087) );
  XNOR2X1_RVT U2832 ( .A1(n1925), .A2(\sub_467/carry[9] ), .Y(N1975) );
  OR2X1_RVT U2833 ( .A1(n1924), .A2(\sub_467/carry[8] ), .Y(\sub_467/carry[9] ) );
  XNOR2X1_RVT U2834 ( .A1(\sub_467/carry[8] ), .A2(n1923), .Y(N1974) );
  OR2X1_RVT U2835 ( .A1(n1922), .A2(\sub_467/carry[7] ), .Y(\sub_467/carry[8] ) );
  XNOR2X1_RVT U2836 ( .A1(\sub_467/carry[7] ), .A2(n1921), .Y(N1973) );
  AND2X1_RVT U2837 ( .A1(n1920), .A2(\sub_467/carry[6] ), .Y(
        \sub_467/carry[7] ) );
  XOR2X1_RVT U2838 ( .A1(n1527), .A2(\sub_467/carry[6] ), .Y(N1972) );
  AND2X1_RVT U2839 ( .A1(n1918), .A2(\sub_467/carry[5] ), .Y(
        \sub_467/carry[6] ) );
  XOR2X1_RVT U2840 ( .A1(n1526), .A2(\sub_467/carry[5] ), .Y(N1971) );
  AND2X1_RVT U2841 ( .A1(n1916), .A2(\sub_467/carry[4] ), .Y(
        \sub_467/carry[5] ) );
  XOR2X1_RVT U2842 ( .A1(n1914), .A2(\sub_467/carry[4] ), .Y(N1970) );
  AND2X1_RVT U2843 ( .A1(n1904), .A2(\sub_467/carry[3] ), .Y(
        \sub_467/carry[4] ) );
  XOR2X1_RVT U2844 ( .A1(n1903), .A2(\sub_467/carry[3] ), .Y(N1969) );
  AND2X1_RVT U2845 ( .A1(n1908), .A2(\sub_467/carry[2] ), .Y(
        \sub_467/carry[3] ) );
  XOR2X1_RVT U2846 ( .A1(n1907), .A2(\sub_467/carry[2] ), .Y(N1968) );
  AND2X1_RVT U2847 ( .A1(n1910), .A2(N1129), .Y(\sub_467/carry[2] ) );
  XOR2X1_RVT U2848 ( .A1(n1909), .A2(N1129), .Y(N1967) );
  XNOR2X1_RVT U2849 ( .A1(n1925), .A2(\sub_368/carry[9] ), .Y(N1533) );
  OR2X1_RVT U2850 ( .A1(n1924), .A2(\sub_368/carry[8] ), .Y(\sub_368/carry[9] ) );
  XNOR2X1_RVT U2851 ( .A1(\sub_368/carry[8] ), .A2(n1923), .Y(N1532) );
  OR2X1_RVT U2852 ( .A1(n1922), .A2(\sub_368/carry[7] ), .Y(\sub_368/carry[8] ) );
  XNOR2X1_RVT U2853 ( .A1(\sub_368/carry[7] ), .A2(n1921), .Y(N1531) );
  OR2X1_RVT U2854 ( .A1(n1920), .A2(\sub_368/carry[6] ), .Y(\sub_368/carry[7] ) );
  XNOR2X1_RVT U2855 ( .A1(\sub_368/carry[6] ), .A2(n1919), .Y(N1530) );
  OR2X1_RVT U2856 ( .A1(n1918), .A2(\sub_368/carry[5] ), .Y(\sub_368/carry[6] ) );
  XNOR2X1_RVT U2857 ( .A1(\sub_368/carry[5] ), .A2(n1917), .Y(N1529) );
  OR2X1_RVT U2858 ( .A1(n1915), .A2(\sub_368/carry[4] ), .Y(\sub_368/carry[5] ) );
  XNOR2X1_RVT U2859 ( .A1(\sub_368/carry[4] ), .A2(n1913), .Y(N1528) );
  AND2X1_RVT U2860 ( .A1(n1904), .A2(\sub_368/carry[3] ), .Y(
        \sub_368/carry[4] ) );
  XOR2X1_RVT U2861 ( .A1(n1903), .A2(\sub_368/carry[3] ), .Y(N1527) );
  OR2X1_RVT U2862 ( .A1(n1908), .A2(\sub_368/carry[2] ), .Y(\sub_368/carry[3] ) );
  XNOR2X1_RVT U2863 ( .A1(\sub_368/carry[2] ), .A2(n1906), .Y(N1526) );
  OR2X1_RVT U2864 ( .A1(n1910), .A2(N1129), .Y(\sub_368/carry[2] ) );
  XNOR2X1_RVT U2865 ( .A1(N1129), .A2(n1909), .Y(N1525) );
  XNOR2X1_RVT U2866 ( .A1(n1925), .A2(\sub_363/carry[9] ), .Y(N1523) );
  OR2X1_RVT U2867 ( .A1(n1924), .A2(\sub_363/carry[8] ), .Y(\sub_363/carry[9] ) );
  XNOR2X1_RVT U2868 ( .A1(\sub_363/carry[8] ), .A2(n1923), .Y(N1522) );
  OR2X1_RVT U2869 ( .A1(n1922), .A2(\sub_363/carry[7] ), .Y(\sub_363/carry[8] ) );
  XNOR2X1_RVT U2870 ( .A1(\sub_363/carry[7] ), .A2(n1921), .Y(N1521) );
  OR2X1_RVT U2871 ( .A1(n1920), .A2(\sub_363/carry[6] ), .Y(\sub_363/carry[7] ) );
  XNOR2X1_RVT U2872 ( .A1(\sub_363/carry[6] ), .A2(n1919), .Y(N1520) );
  OR2X1_RVT U2873 ( .A1(n1918), .A2(\sub_363/carry[5] ), .Y(\sub_363/carry[6] ) );
  XNOR2X1_RVT U2874 ( .A1(\sub_363/carry[5] ), .A2(n1917), .Y(N1519) );
  OR2X1_RVT U2875 ( .A1(n1915), .A2(\sub_363/carry[4] ), .Y(\sub_363/carry[5] ) );
  XNOR2X1_RVT U2876 ( .A1(\sub_363/carry[4] ), .A2(n1913), .Y(N1518) );
  AND2X1_RVT U2877 ( .A1(n1904), .A2(\sub_363/carry[3] ), .Y(
        \sub_363/carry[4] ) );
  XOR2X1_RVT U2878 ( .A1(n1903), .A2(\sub_363/carry[3] ), .Y(N1517) );
  OR2X1_RVT U2879 ( .A1(n1908), .A2(n1909), .Y(\sub_363/carry[3] ) );
  XNOR2X1_RVT U2880 ( .A1(n1909), .A2(n1906), .Y(N1516) );
  XNOR2X1_RVT U2881 ( .A1(n1925), .A2(\sub_304/carry[9] ), .Y(N1266) );
  OR2X1_RVT U2882 ( .A1(n1924), .A2(\sub_304/carry[8] ), .Y(\sub_304/carry[9] ) );
  XNOR2X1_RVT U2883 ( .A1(\sub_304/carry[8] ), .A2(n1923), .Y(N1265) );
  OR2X1_RVT U2884 ( .A1(n1922), .A2(\sub_304/carry[7] ), .Y(\sub_304/carry[8] ) );
  XNOR2X1_RVT U2885 ( .A1(\sub_304/carry[7] ), .A2(n1921), .Y(N1264) );
  OR2X1_RVT U2886 ( .A1(n1920), .A2(\sub_304/carry[6] ), .Y(\sub_304/carry[7] ) );
  XNOR2X1_RVT U2887 ( .A1(\sub_304/carry[6] ), .A2(n1919), .Y(N1263) );
  OR2X1_RVT U2888 ( .A1(n1918), .A2(\sub_304/carry[5] ), .Y(\sub_304/carry[6] ) );
  XNOR2X1_RVT U2889 ( .A1(\sub_304/carry[5] ), .A2(n1917), .Y(N1262) );
  AND2X1_RVT U2890 ( .A1(n1915), .A2(\sub_304/carry[4] ), .Y(
        \sub_304/carry[5] ) );
  XOR2X1_RVT U2891 ( .A1(n1914), .A2(\sub_304/carry[4] ), .Y(N1261) );
  OR2X1_RVT U2892 ( .A1(n1904), .A2(\sub_304/carry[3] ), .Y(\sub_304/carry[4] ) );
  XNOR2X1_RVT U2893 ( .A1(\sub_304/carry[3] ), .A2(n1902), .Y(N1260) );
  OR2X1_RVT U2894 ( .A1(n1908), .A2(\sub_304/carry[2] ), .Y(\sub_304/carry[3] ) );
  XNOR2X1_RVT U2895 ( .A1(\sub_304/carry[2] ), .A2(n1906), .Y(N1259) );
  OR2X1_RVT U2896 ( .A1(n1909), .A2(N1129), .Y(\sub_304/carry[2] ) );
  XNOR2X1_RVT U2897 ( .A1(N1129), .A2(n1909), .Y(N1258) );
  XNOR2X1_RVT U2898 ( .A1(n1925), .A2(\sub_299/carry[9] ), .Y(N1256) );
  OR2X1_RVT U2899 ( .A1(n1924), .A2(\sub_299/carry[8] ), .Y(\sub_299/carry[9] ) );
  XNOR2X1_RVT U2900 ( .A1(\sub_299/carry[8] ), .A2(n1923), .Y(N1255) );
  OR2X1_RVT U2901 ( .A1(n1922), .A2(\sub_299/carry[7] ), .Y(\sub_299/carry[8] ) );
  XNOR2X1_RVT U2902 ( .A1(\sub_299/carry[7] ), .A2(n1921), .Y(N1254) );
  OR2X1_RVT U2903 ( .A1(n1920), .A2(\sub_299/carry[6] ), .Y(\sub_299/carry[7] ) );
  XNOR2X1_RVT U2904 ( .A1(\sub_299/carry[6] ), .A2(n1919), .Y(N1253) );
  OR2X1_RVT U2905 ( .A1(n1918), .A2(\sub_299/carry[5] ), .Y(\sub_299/carry[6] ) );
  XNOR2X1_RVT U2906 ( .A1(\sub_299/carry[5] ), .A2(n1917), .Y(N1252) );
  AND2X1_RVT U2907 ( .A1(n1915), .A2(\sub_299/carry[4] ), .Y(
        \sub_299/carry[5] ) );
  XOR2X1_RVT U2908 ( .A1(n1914), .A2(\sub_299/carry[4] ), .Y(N1251) );
  OR2X1_RVT U2909 ( .A1(n1904), .A2(\sub_299/carry[3] ), .Y(\sub_299/carry[4] ) );
  XNOR2X1_RVT U2910 ( .A1(\sub_299/carry[3] ), .A2(n1902), .Y(N1250) );
  OR2X1_RVT U2911 ( .A1(n1908), .A2(n1909), .Y(\sub_299/carry[3] ) );
  XNOR2X1_RVT U2912 ( .A1(n1909), .A2(n1906), .Y(N1249) );
  XNOR2X1_RVT U2913 ( .A1(n1925), .A2(\sub_288/carry[9] ), .Y(N1206) );
  OR2X1_RVT U2914 ( .A1(n1924), .A2(\sub_288/carry[8] ), .Y(\sub_288/carry[9] ) );
  XNOR2X1_RVT U2915 ( .A1(\sub_288/carry[8] ), .A2(n1923), .Y(N1205) );
  OR2X1_RVT U2916 ( .A1(n1922), .A2(\sub_288/carry[7] ), .Y(\sub_288/carry[8] ) );
  XNOR2X1_RVT U2917 ( .A1(\sub_288/carry[7] ), .A2(n1921), .Y(N1204) );
  OR2X1_RVT U2918 ( .A1(n1920), .A2(\sub_288/carry[6] ), .Y(\sub_288/carry[7] ) );
  XNOR2X1_RVT U2919 ( .A1(\sub_288/carry[6] ), .A2(n1919), .Y(N1203) );
  OR2X1_RVT U2920 ( .A1(n1918), .A2(\sub_288/carry[5] ), .Y(\sub_288/carry[6] ) );
  XNOR2X1_RVT U2921 ( .A1(\sub_288/carry[5] ), .A2(n1917), .Y(N1202) );
  AND2X1_RVT U2922 ( .A1(n1915), .A2(\sub_288/carry[4] ), .Y(
        \sub_288/carry[5] ) );
  XOR2X1_RVT U2923 ( .A1(n1914), .A2(\sub_288/carry[4] ), .Y(N1201) );
  OR2X1_RVT U2924 ( .A1(n1904), .A2(\sub_288/carry[3] ), .Y(\sub_288/carry[4] ) );
  XNOR2X1_RVT U2925 ( .A1(\sub_288/carry[3] ), .A2(n1902), .Y(N1200) );
  OR2X1_RVT U2926 ( .A1(n1908), .A2(\sub_288/carry[2] ), .Y(\sub_288/carry[3] ) );
  XNOR2X1_RVT U2927 ( .A1(\sub_288/carry[2] ), .A2(n1906), .Y(N1199) );
  AND2X1_RVT U2928 ( .A1(n1910), .A2(N1129), .Y(\sub_288/carry[2] ) );
  XOR2X1_RVT U2929 ( .A1(n1909), .A2(N1129), .Y(N1198) );
  XNOR2X1_RVT U2930 ( .A1(n1925), .A2(\sub_352/carry[9] ), .Y(N1465) );
  OR2X1_RVT U2931 ( .A1(n1924), .A2(\sub_352/carry[8] ), .Y(\sub_352/carry[9] ) );
  XNOR2X1_RVT U2932 ( .A1(\sub_352/carry[8] ), .A2(n1923), .Y(N1464) );
  OR2X1_RVT U2933 ( .A1(n1922), .A2(\sub_352/carry[7] ), .Y(\sub_352/carry[8] ) );
  XNOR2X1_RVT U2934 ( .A1(\sub_352/carry[7] ), .A2(n1921), .Y(N1463) );
  OR2X1_RVT U2935 ( .A1(n1920), .A2(\sub_352/carry[6] ), .Y(\sub_352/carry[7] ) );
  XNOR2X1_RVT U2936 ( .A1(\sub_352/carry[6] ), .A2(n1919), .Y(N1462) );
  OR2X1_RVT U2937 ( .A1(n1918), .A2(\sub_352/carry[5] ), .Y(\sub_352/carry[6] ) );
  XNOR2X1_RVT U2938 ( .A1(\sub_352/carry[5] ), .A2(n1917), .Y(N1461) );
  OR2X1_RVT U2939 ( .A1(n1915), .A2(\sub_352/carry[4] ), .Y(\sub_352/carry[5] ) );
  XNOR2X1_RVT U2940 ( .A1(\sub_352/carry[4] ), .A2(n1913), .Y(N1460) );
  AND2X1_RVT U2941 ( .A1(n1904), .A2(\sub_352/carry[3] ), .Y(
        \sub_352/carry[4] ) );
  XOR2X1_RVT U2942 ( .A1(n1903), .A2(\sub_352/carry[3] ), .Y(N1459) );
  OR2X1_RVT U2943 ( .A1(n1908), .A2(\sub_352/carry[2] ), .Y(\sub_352/carry[3] ) );
  XNOR2X1_RVT U2944 ( .A1(\sub_352/carry[2] ), .A2(n1906), .Y(N1458) );
  AND2X1_RVT U2945 ( .A1(n1910), .A2(N1129), .Y(\sub_352/carry[2] ) );
  XOR2X1_RVT U2946 ( .A1(n1909), .A2(N1129), .Y(N1457) );
  XNOR2X1_RVT U2947 ( .A1(n1925), .A2(\sub_347/carry[9] ), .Y(N1455) );
  OR2X1_RVT U2948 ( .A1(n1924), .A2(\sub_347/carry[8] ), .Y(\sub_347/carry[9] ) );
  XNOR2X1_RVT U2949 ( .A1(\sub_347/carry[8] ), .A2(n1923), .Y(N1454) );
  OR2X1_RVT U2950 ( .A1(n1922), .A2(\sub_347/carry[7] ), .Y(\sub_347/carry[8] ) );
  XNOR2X1_RVT U2951 ( .A1(\sub_347/carry[7] ), .A2(n1921), .Y(N1453) );
  OR2X1_RVT U2952 ( .A1(n1920), .A2(\sub_347/carry[6] ), .Y(\sub_347/carry[7] ) );
  XNOR2X1_RVT U2953 ( .A1(\sub_347/carry[6] ), .A2(n1919), .Y(N1452) );
  OR2X1_RVT U2954 ( .A1(n1918), .A2(\sub_347/carry[5] ), .Y(\sub_347/carry[6] ) );
  XNOR2X1_RVT U2955 ( .A1(\sub_347/carry[5] ), .A2(n1917), .Y(N1451) );
  OR2X1_RVT U2956 ( .A1(n1915), .A2(\sub_347/carry[4] ), .Y(\sub_347/carry[5] ) );
  XNOR2X1_RVT U2957 ( .A1(\sub_347/carry[4] ), .A2(n1913), .Y(N1450) );
  AND2X1_RVT U2958 ( .A1(n1904), .A2(n1908), .Y(\sub_347/carry[4] ) );
  XOR2X1_RVT U2959 ( .A1(n1903), .A2(n1906), .Y(N1449) );
  XNOR2X1_RVT U2960 ( .A1(n1925), .A2(\sub_339/carry[9] ), .Y(N1399) );
  OR2X1_RVT U2961 ( .A1(n1924), .A2(\sub_339/carry[8] ), .Y(\sub_339/carry[9] ) );
  XNOR2X1_RVT U2962 ( .A1(\sub_339/carry[8] ), .A2(n1923), .Y(N1398) );
  OR2X1_RVT U2963 ( .A1(n1922), .A2(\sub_339/carry[7] ), .Y(\sub_339/carry[8] ) );
  XNOR2X1_RVT U2964 ( .A1(\sub_339/carry[7] ), .A2(n1921), .Y(N1397) );
  OR2X1_RVT U2965 ( .A1(n1920), .A2(\sub_339/carry[6] ), .Y(\sub_339/carry[7] ) );
  XNOR2X1_RVT U2966 ( .A1(\sub_339/carry[6] ), .A2(n1919), .Y(N1396) );
  OR2X1_RVT U2967 ( .A1(n1918), .A2(\sub_339/carry[5] ), .Y(\sub_339/carry[6] ) );
  XNOR2X1_RVT U2968 ( .A1(\sub_339/carry[5] ), .A2(n1917), .Y(N1395) );
  OR2X1_RVT U2969 ( .A1(n1915), .A2(\sub_339/carry[4] ), .Y(\sub_339/carry[5] ) );
  XNOR2X1_RVT U2970 ( .A1(\sub_339/carry[4] ), .A2(n1914), .Y(N1394) );
  AND2X1_RVT U2971 ( .A1(n1904), .A2(\sub_339/carry[3] ), .Y(
        \sub_339/carry[4] ) );
  XOR2X1_RVT U2972 ( .A1(n1903), .A2(\sub_339/carry[3] ), .Y(N1393) );
  AND2X1_RVT U2973 ( .A1(n1908), .A2(\sub_339/carry[2] ), .Y(
        \sub_339/carry[3] ) );
  XOR2X1_RVT U2974 ( .A1(n1907), .A2(\sub_339/carry[2] ), .Y(N1392) );
  OR2X1_RVT U2975 ( .A1(n1910), .A2(N1129), .Y(\sub_339/carry[2] ) );
  XNOR2X1_RVT U2976 ( .A1(N1129), .A2(n1909), .Y(N1391) );
  XNOR2X1_RVT U2977 ( .A1(n1925), .A2(\sub_283/carry[9] ), .Y(N1196) );
  OR2X1_RVT U2978 ( .A1(n1924), .A2(\sub_283/carry[8] ), .Y(\sub_283/carry[9] ) );
  XNOR2X1_RVT U2979 ( .A1(\sub_283/carry[8] ), .A2(n1528), .Y(N1195) );
  OR2X1_RVT U2980 ( .A1(n1922), .A2(\sub_283/carry[7] ), .Y(\sub_283/carry[8] ) );
  XNOR2X1_RVT U2981 ( .A1(\sub_283/carry[7] ), .A2(n1525), .Y(N1194) );
  OR2X1_RVT U2982 ( .A1(n1920), .A2(\sub_283/carry[6] ), .Y(\sub_283/carry[7] ) );
  XNOR2X1_RVT U2983 ( .A1(\sub_283/carry[6] ), .A2(n1527), .Y(N1193) );
  OR2X1_RVT U2984 ( .A1(n1918), .A2(\sub_283/carry[5] ), .Y(\sub_283/carry[6] ) );
  XNOR2X1_RVT U2985 ( .A1(\sub_283/carry[5] ), .A2(n1526), .Y(N1192) );
  AND2X1_RVT U2986 ( .A1(n1915), .A2(\sub_283/carry[4] ), .Y(
        \sub_283/carry[5] ) );
  XOR2X1_RVT U2987 ( .A1(n1914), .A2(\sub_283/carry[4] ), .Y(N1191) );
  OR2X1_RVT U2988 ( .A1(n1904), .A2(n1907), .Y(\sub_283/carry[4] ) );
  XNOR2X1_RVT U2989 ( .A1(n1906), .A2(n1902), .Y(N1190) );
  XNOR2X1_RVT U2990 ( .A1(n1925), .A2(\sub_270/carry[9] ), .Y(N1138) );
  OR2X1_RVT U2991 ( .A1(n1924), .A2(\sub_270/carry[8] ), .Y(\sub_270/carry[9] ) );
  XNOR2X1_RVT U2992 ( .A1(\sub_270/carry[8] ), .A2(n1528), .Y(N1137) );
  OR2X1_RVT U2993 ( .A1(n1922), .A2(\sub_270/carry[7] ), .Y(\sub_270/carry[8] ) );
  XNOR2X1_RVT U2994 ( .A1(\sub_270/carry[7] ), .A2(n1921), .Y(N1136) );
  OR2X1_RVT U2995 ( .A1(n1920), .A2(\sub_270/carry[6] ), .Y(\sub_270/carry[7] ) );
  XNOR2X1_RVT U2996 ( .A1(\sub_270/carry[6] ), .A2(n1919), .Y(N1135) );
  OR2X1_RVT U2997 ( .A1(n1918), .A2(\sub_270/carry[5] ), .Y(\sub_270/carry[6] ) );
  XNOR2X1_RVT U2998 ( .A1(\sub_270/carry[5] ), .A2(n1917), .Y(N1134) );
  AND2X1_RVT U2999 ( .A1(n1915), .A2(\sub_270/carry[4] ), .Y(
        \sub_270/carry[5] ) );
  XOR2X1_RVT U3000 ( .A1(n1914), .A2(\sub_270/carry[4] ), .Y(N1133) );
  OR2X1_RVT U3001 ( .A1(n1904), .A2(\sub_270/carry[3] ), .Y(\sub_270/carry[4] ) );
  XNOR2X1_RVT U3002 ( .A1(\sub_270/carry[3] ), .A2(n1902), .Y(N1132) );
  AND2X1_RVT U3003 ( .A1(n1908), .A2(n1910), .Y(\sub_270/carry[3] ) );
  XOR2X1_RVT U3004 ( .A1(n1907), .A2(n1909), .Y(N1131) );
  XNOR2X1_RVT U3005 ( .A1(n1925), .A2(\sub_259/carry[9] ), .Y(N1124) );
  OR2X1_RVT U3006 ( .A1(n1924), .A2(\sub_259/carry[8] ), .Y(\sub_259/carry[9] ) );
  XNOR2X1_RVT U3007 ( .A1(\sub_259/carry[8] ), .A2(n1528), .Y(N1123) );
  OR2X1_RVT U3008 ( .A1(n1922), .A2(\sub_259/carry[7] ), .Y(\sub_259/carry[8] ) );
  XNOR2X1_RVT U3009 ( .A1(\sub_259/carry[7] ), .A2(n1921), .Y(N1122) );
  OR2X1_RVT U3010 ( .A1(n1920), .A2(\sub_259/carry[6] ), .Y(\sub_259/carry[7] ) );
  XNOR2X1_RVT U3011 ( .A1(\sub_259/carry[6] ), .A2(n1919), .Y(N1121) );
  OR2X1_RVT U3012 ( .A1(n1918), .A2(\sub_259/carry[5] ), .Y(\sub_259/carry[6] ) );
  XNOR2X1_RVT U3013 ( .A1(\sub_259/carry[5] ), .A2(n1917), .Y(N1120) );
  AND2X1_RVT U3014 ( .A1(n1915), .A2(\sub_259/carry[4] ), .Y(
        \sub_259/carry[5] ) );
  XOR2X1_RVT U3015 ( .A1(n1914), .A2(\sub_259/carry[4] ), .Y(N1119) );
  OR2X1_RVT U3016 ( .A1(n1904), .A2(\sub_259/carry[3] ), .Y(\sub_259/carry[4] ) );
  XNOR2X1_RVT U3017 ( .A1(\sub_259/carry[3] ), .A2(n1903), .Y(N1118) );
  AND2X1_RVT U3018 ( .A1(n1908), .A2(\sub_259/carry[2] ), .Y(
        \sub_259/carry[3] ) );
  XOR2X1_RVT U3019 ( .A1(n1907), .A2(\sub_259/carry[2] ), .Y(N1117) );
  AND2X1_RVT U3020 ( .A1(n1910), .A2(N1129), .Y(\sub_259/carry[2] ) );
  XOR2X1_RVT U3021 ( .A1(n1909), .A2(N1129), .Y(N1116) );
  XNOR2X1_RVT U3022 ( .A1(n1926), .A2(\sub_275/carry[9] ), .Y(N1148) );
  OR2X1_RVT U3023 ( .A1(n1924), .A2(\sub_275/carry[8] ), .Y(\sub_275/carry[9] ) );
  XNOR2X1_RVT U3024 ( .A1(\sub_275/carry[8] ), .A2(n1528), .Y(N1147) );
  OR2X1_RVT U3025 ( .A1(n1922), .A2(\sub_275/carry[7] ), .Y(\sub_275/carry[8] ) );
  XNOR2X1_RVT U3026 ( .A1(\sub_275/carry[7] ), .A2(n1921), .Y(N1146) );
  OR2X1_RVT U3027 ( .A1(n1920), .A2(\sub_275/carry[6] ), .Y(\sub_275/carry[7] ) );
  XNOR2X1_RVT U3028 ( .A1(\sub_275/carry[6] ), .A2(n1919), .Y(N1145) );
  OR2X1_RVT U3029 ( .A1(n1918), .A2(\sub_275/carry[5] ), .Y(\sub_275/carry[6] ) );
  XNOR2X1_RVT U3030 ( .A1(\sub_275/carry[5] ), .A2(n1917), .Y(N1144) );
  AND2X1_RVT U3031 ( .A1(n1915), .A2(\sub_275/carry[4] ), .Y(
        \sub_275/carry[5] ) );
  XOR2X1_RVT U3032 ( .A1(n1914), .A2(\sub_275/carry[4] ), .Y(N1143) );
  OR2X1_RVT U3033 ( .A1(n1904), .A2(\sub_275/carry[3] ), .Y(\sub_275/carry[4] ) );
  XNOR2X1_RVT U3034 ( .A1(\sub_275/carry[3] ), .A2(n1903), .Y(N1142) );
  AND2X1_RVT U3035 ( .A1(n1908), .A2(\sub_275/carry[2] ), .Y(
        \sub_275/carry[3] ) );
  XOR2X1_RVT U3036 ( .A1(n1907), .A2(\sub_275/carry[2] ), .Y(N1141) );
  OR2X1_RVT U3037 ( .A1(n1909), .A2(N1129), .Y(\sub_275/carry[2] ) );
  XNOR2X1_RVT U3038 ( .A1(N1129), .A2(n1909), .Y(N1140) );
  XNOR2X1_RVT U3039 ( .A1(n1926), .A2(\sub_334/carry[9] ), .Y(N1389) );
  OR2X1_RVT U3040 ( .A1(n1924), .A2(\sub_334/carry[8] ), .Y(\sub_334/carry[9] ) );
  XNOR2X1_RVT U3041 ( .A1(\sub_334/carry[8] ), .A2(n1528), .Y(N1388) );
  OR2X1_RVT U3042 ( .A1(n1922), .A2(\sub_334/carry[7] ), .Y(\sub_334/carry[8] ) );
  XNOR2X1_RVT U3043 ( .A1(\sub_334/carry[7] ), .A2(n1921), .Y(N1387) );
  OR2X1_RVT U3044 ( .A1(n1920), .A2(\sub_334/carry[6] ), .Y(\sub_334/carry[7] ) );
  XNOR2X1_RVT U3045 ( .A1(\sub_334/carry[6] ), .A2(n1919), .Y(N1386) );
  OR2X1_RVT U3046 ( .A1(n1918), .A2(\sub_334/carry[5] ), .Y(\sub_334/carry[6] ) );
  XNOR2X1_RVT U3047 ( .A1(\sub_334/carry[5] ), .A2(n1917), .Y(N1385) );
  OR2X1_RVT U3048 ( .A1(n1915), .A2(\sub_334/carry[4] ), .Y(\sub_334/carry[5] ) );
  XNOR2X1_RVT U3049 ( .A1(\sub_334/carry[4] ), .A2(n1914), .Y(N1384) );
  AND2X1_RVT U3050 ( .A1(n1904), .A2(\sub_334/carry[3] ), .Y(
        \sub_334/carry[4] ) );
  XOR2X1_RVT U3051 ( .A1(n1903), .A2(\sub_334/carry[3] ), .Y(N1383) );
  AND2X1_RVT U3052 ( .A1(n1908), .A2(n1910), .Y(\sub_334/carry[3] ) );
  XOR2X1_RVT U3053 ( .A1(n1907), .A2(n1909), .Y(N1382) );
  XNOR2X1_RVT U3054 ( .A1(n1926), .A2(\sub_400/carry[9] ), .Y(N1678) );
  OR2X1_RVT U3055 ( .A1(n1924), .A2(\sub_400/carry[8] ), .Y(\sub_400/carry[9] ) );
  XNOR2X1_RVT U3056 ( .A1(\sub_400/carry[8] ), .A2(n1528), .Y(N1677) );
  OR2X1_RVT U3057 ( .A1(n1922), .A2(\sub_400/carry[7] ), .Y(\sub_400/carry[8] ) );
  XNOR2X1_RVT U3058 ( .A1(\sub_400/carry[7] ), .A2(n1921), .Y(N1676) );
  OR2X1_RVT U3059 ( .A1(n1920), .A2(\sub_400/carry[6] ), .Y(\sub_400/carry[7] ) );
  XNOR2X1_RVT U3060 ( .A1(\sub_400/carry[6] ), .A2(n1919), .Y(N1675) );
  OR2X1_RVT U3061 ( .A1(n1918), .A2(\sub_400/carry[5] ), .Y(\sub_400/carry[6] ) );
  XNOR2X1_RVT U3062 ( .A1(\sub_400/carry[5] ), .A2(n1917), .Y(N1674) );
  OR2X1_RVT U3063 ( .A1(n1915), .A2(\sub_400/carry[4] ), .Y(\sub_400/carry[5] ) );
  XNOR2X1_RVT U3064 ( .A1(\sub_400/carry[4] ), .A2(n1914), .Y(N1673) );
  OR2X1_RVT U3065 ( .A1(n1904), .A2(\sub_400/carry[3] ), .Y(\sub_400/carry[4] ) );
  XNOR2X1_RVT U3066 ( .A1(\sub_400/carry[3] ), .A2(n1903), .Y(N1672) );
  AND2X1_RVT U3067 ( .A1(n1908), .A2(\sub_400/carry[2] ), .Y(
        \sub_400/carry[3] ) );
  XOR2X1_RVT U3068 ( .A1(n1907), .A2(\sub_400/carry[2] ), .Y(N1671) );
  OR2X1_RVT U3069 ( .A1(n1909), .A2(n1911), .Y(\sub_400/carry[2] ) );
  XNOR2X1_RVT U3070 ( .A1(N1129), .A2(n1909), .Y(N1670) );
  XNOR2X1_RVT U3071 ( .A1(n1926), .A2(\sub_424/carry[9] ), .Y(N1818) );
  OR2X1_RVT U3072 ( .A1(n1924), .A2(\sub_424/carry[8] ), .Y(\sub_424/carry[9] ) );
  XNOR2X1_RVT U3073 ( .A1(\sub_424/carry[8] ), .A2(n1923), .Y(N1817) );
  OR2X1_RVT U3074 ( .A1(n1525), .A2(\sub_424/carry[7] ), .Y(\sub_424/carry[8] ) );
  XNOR2X1_RVT U3075 ( .A1(\sub_424/carry[7] ), .A2(n1525), .Y(N1816) );
  OR2X1_RVT U3076 ( .A1(n1527), .A2(\sub_424/carry[6] ), .Y(\sub_424/carry[7] ) );
  XNOR2X1_RVT U3077 ( .A1(\sub_424/carry[6] ), .A2(n1919), .Y(N1815) );
  OR2X1_RVT U3078 ( .A1(n1526), .A2(\sub_424/carry[5] ), .Y(\sub_424/carry[6] ) );
  XNOR2X1_RVT U3079 ( .A1(\sub_424/carry[5] ), .A2(n1917), .Y(N1814) );
  OR2X1_RVT U3080 ( .A1(n1915), .A2(\sub_424/carry[4] ), .Y(\sub_424/carry[5] ) );
  XNOR2X1_RVT U3081 ( .A1(\sub_424/carry[4] ), .A2(n1914), .Y(N1813) );
  OR2X1_RVT U3082 ( .A1(n1904), .A2(\sub_424/carry[3] ), .Y(\sub_424/carry[4] ) );
  XNOR2X1_RVT U3083 ( .A1(\sub_424/carry[3] ), .A2(n1902), .Y(N1812) );
  OR2X1_RVT U3084 ( .A1(n1908), .A2(n1909), .Y(\sub_424/carry[3] ) );
  XNOR2X1_RVT U3085 ( .A1(n1909), .A2(n1906), .Y(N1811) );
  XNOR2X1_RVT U3086 ( .A1(n1926), .A2(\sub_395/carry[9] ), .Y(N1668) );
  OR2X1_RVT U3087 ( .A1(n1924), .A2(\sub_395/carry[8] ), .Y(\sub_395/carry[9] ) );
  XNOR2X1_RVT U3088 ( .A1(\sub_395/carry[8] ), .A2(n1528), .Y(N1667) );
  OR2X1_RVT U3089 ( .A1(n1525), .A2(\sub_395/carry[7] ), .Y(\sub_395/carry[8] ) );
  XNOR2X1_RVT U3090 ( .A1(\sub_395/carry[7] ), .A2(n1525), .Y(N1666) );
  OR2X1_RVT U3091 ( .A1(n1527), .A2(\sub_395/carry[6] ), .Y(\sub_395/carry[7] ) );
  XNOR2X1_RVT U3092 ( .A1(\sub_395/carry[6] ), .A2(n1527), .Y(N1665) );
  OR2X1_RVT U3093 ( .A1(n1526), .A2(\sub_395/carry[5] ), .Y(\sub_395/carry[6] ) );
  XNOR2X1_RVT U3094 ( .A1(\sub_395/carry[5] ), .A2(n1526), .Y(N1664) );
  OR2X1_RVT U3095 ( .A1(n1915), .A2(\sub_395/carry[4] ), .Y(\sub_395/carry[5] ) );
  XNOR2X1_RVT U3096 ( .A1(\sub_395/carry[4] ), .A2(n1913), .Y(N1663) );
  OR2X1_RVT U3097 ( .A1(n1904), .A2(\sub_395/carry[3] ), .Y(\sub_395/carry[4] ) );
  XNOR2X1_RVT U3098 ( .A1(\sub_395/carry[3] ), .A2(n1902), .Y(N1662) );
  AND2X1_RVT U3099 ( .A1(n1908), .A2(n1910), .Y(\sub_395/carry[3] ) );
  XOR2X1_RVT U3100 ( .A1(n1907), .A2(n1909), .Y(N1661) );
  XNOR2X1_RVT U3101 ( .A1(n1926), .A2(\sub_408/carry[9] ), .Y(N1742) );
  OR2X1_RVT U3102 ( .A1(n1924), .A2(\sub_408/carry[8] ), .Y(\sub_408/carry[9] ) );
  XNOR2X1_RVT U3103 ( .A1(\sub_408/carry[8] ), .A2(n1528), .Y(N1741) );
  OR2X1_RVT U3104 ( .A1(n1922), .A2(\sub_408/carry[7] ), .Y(\sub_408/carry[8] ) );
  XNOR2X1_RVT U3105 ( .A1(\sub_408/carry[7] ), .A2(n1525), .Y(N1740) );
  OR2X1_RVT U3106 ( .A1(n1920), .A2(\sub_408/carry[6] ), .Y(\sub_408/carry[7] ) );
  XNOR2X1_RVT U3107 ( .A1(\sub_408/carry[6] ), .A2(n1527), .Y(N1739) );
  OR2X1_RVT U3108 ( .A1(n1918), .A2(\sub_408/carry[5] ), .Y(\sub_408/carry[6] ) );
  XNOR2X1_RVT U3109 ( .A1(\sub_408/carry[5] ), .A2(n1526), .Y(N1738) );
  OR2X1_RVT U3110 ( .A1(n1915), .A2(\sub_408/carry[4] ), .Y(\sub_408/carry[5] ) );
  XNOR2X1_RVT U3111 ( .A1(\sub_408/carry[4] ), .A2(n1913), .Y(N1737) );
  OR2X1_RVT U3112 ( .A1(n1904), .A2(n1907), .Y(\sub_408/carry[4] ) );
  XNOR2X1_RVT U3113 ( .A1(n1906), .A2(n1902), .Y(N1736) );
  XNOR2X1_RVT U3114 ( .A1(n1926), .A2(\sub_317/carry[9] ), .Y(N1328) );
  OR2X1_RVT U3115 ( .A1(n1528), .A2(\sub_317/carry[8] ), .Y(\sub_317/carry[9] ) );
  XNOR2X1_RVT U3116 ( .A1(\sub_317/carry[8] ), .A2(n1528), .Y(N1327) );
  OR2X1_RVT U3117 ( .A1(n1922), .A2(\sub_317/carry[7] ), .Y(\sub_317/carry[8] ) );
  XNOR2X1_RVT U3118 ( .A1(\sub_317/carry[7] ), .A2(n1525), .Y(N1326) );
  OR2X1_RVT U3119 ( .A1(n1527), .A2(\sub_317/carry[6] ), .Y(\sub_317/carry[7] ) );
  XNOR2X1_RVT U3120 ( .A1(\sub_317/carry[6] ), .A2(n1527), .Y(N1325) );
  OR2X1_RVT U3121 ( .A1(n1526), .A2(\sub_317/carry[5] ), .Y(\sub_317/carry[6] ) );
  XNOR2X1_RVT U3122 ( .A1(\sub_317/carry[5] ), .A2(n1526), .Y(N1324) );
  OR2X1_RVT U3123 ( .A1(n1915), .A2(\sub_317/carry[4] ), .Y(\sub_317/carry[5] ) );
  XNOR2X1_RVT U3124 ( .A1(\sub_317/carry[4] ), .A2(n1913), .Y(N1323) );
  AND2X1_RVT U3125 ( .A1(n1904), .A2(\sub_317/carry[3] ), .Y(
        \sub_317/carry[4] ) );
  XOR2X1_RVT U3126 ( .A1(n1903), .A2(\sub_317/carry[3] ), .Y(N1322) );
  AND2X1_RVT U3127 ( .A1(n1908), .A2(\sub_317/carry[2] ), .Y(
        \sub_317/carry[3] ) );
  XOR2X1_RVT U3128 ( .A1(n1907), .A2(\sub_317/carry[2] ), .Y(N1321) );
  AND2X1_RVT U3129 ( .A1(n1910), .A2(N1129), .Y(\sub_317/carry[2] ) );
  XOR2X1_RVT U3130 ( .A1(n1909), .A2(N1129), .Y(N1320) );
  XNOR2X1_RVT U3131 ( .A1(n1926), .A2(\sub_413/carry[9] ), .Y(N1752) );
  OR2X1_RVT U3132 ( .A1(n1528), .A2(\sub_413/carry[8] ), .Y(\sub_413/carry[9] ) );
  XNOR2X1_RVT U3133 ( .A1(\sub_413/carry[8] ), .A2(n1528), .Y(N1751) );
  OR2X1_RVT U3134 ( .A1(n1525), .A2(\sub_413/carry[7] ), .Y(\sub_413/carry[8] ) );
  XNOR2X1_RVT U3135 ( .A1(\sub_413/carry[7] ), .A2(n1525), .Y(N1750) );
  OR2X1_RVT U3136 ( .A1(n1920), .A2(\sub_413/carry[6] ), .Y(\sub_413/carry[7] ) );
  XNOR2X1_RVT U3137 ( .A1(\sub_413/carry[6] ), .A2(n1527), .Y(N1749) );
  OR2X1_RVT U3138 ( .A1(n1918), .A2(\sub_413/carry[5] ), .Y(\sub_413/carry[6] ) );
  XNOR2X1_RVT U3139 ( .A1(\sub_413/carry[5] ), .A2(n1526), .Y(N1748) );
  OR2X1_RVT U3140 ( .A1(n1915), .A2(\sub_413/carry[4] ), .Y(\sub_413/carry[5] ) );
  XNOR2X1_RVT U3141 ( .A1(\sub_413/carry[4] ), .A2(n1913), .Y(N1747) );
  OR2X1_RVT U3142 ( .A1(n1904), .A2(\sub_413/carry[3] ), .Y(\sub_413/carry[4] ) );
  XNOR2X1_RVT U3143 ( .A1(\sub_413/carry[3] ), .A2(n1902), .Y(N1746) );
  OR2X1_RVT U3144 ( .A1(n1907), .A2(\sub_413/carry[2] ), .Y(\sub_413/carry[3] ) );
  XNOR2X1_RVT U3145 ( .A1(\sub_413/carry[2] ), .A2(n1906), .Y(N1745) );
  AND2X1_RVT U3146 ( .A1(n1910), .A2(N1129), .Y(\sub_413/carry[2] ) );
  XOR2X1_RVT U3147 ( .A1(n1909), .A2(N1129), .Y(N1744) );
  XNOR2X1_RVT U3148 ( .A1(n1926), .A2(\sub_381/carry[9] ), .Y(N1603) );
  OR2X1_RVT U3149 ( .A1(n1924), .A2(\sub_381/carry[8] ), .Y(\sub_381/carry[9] ) );
  XNOR2X1_RVT U3150 ( .A1(\sub_381/carry[8] ), .A2(n1923), .Y(N1602) );
  OR2X1_RVT U3151 ( .A1(n1922), .A2(\sub_381/carry[7] ), .Y(\sub_381/carry[8] ) );
  XNOR2X1_RVT U3152 ( .A1(\sub_381/carry[7] ), .A2(n1525), .Y(N1601) );
  OR2X1_RVT U3153 ( .A1(n1920), .A2(\sub_381/carry[6] ), .Y(\sub_381/carry[7] ) );
  XNOR2X1_RVT U3154 ( .A1(\sub_381/carry[6] ), .A2(n1527), .Y(N1600) );
  OR2X1_RVT U3155 ( .A1(n1918), .A2(\sub_381/carry[5] ), .Y(\sub_381/carry[6] ) );
  XNOR2X1_RVT U3156 ( .A1(\sub_381/carry[5] ), .A2(n1526), .Y(N1599) );
  OR2X1_RVT U3157 ( .A1(n1915), .A2(\sub_381/carry[4] ), .Y(\sub_381/carry[5] ) );
  XNOR2X1_RVT U3158 ( .A1(\sub_381/carry[4] ), .A2(n1913), .Y(N1598) );
  OR2X1_RVT U3159 ( .A1(n1904), .A2(\sub_381/carry[3] ), .Y(\sub_381/carry[4] ) );
  XNOR2X1_RVT U3160 ( .A1(\sub_381/carry[3] ), .A2(n1902), .Y(N1597) );
  AND2X1_RVT U3161 ( .A1(n1908), .A2(\sub_381/carry[2] ), .Y(
        \sub_381/carry[3] ) );
  XOR2X1_RVT U3162 ( .A1(n1907), .A2(\sub_381/carry[2] ), .Y(N1596) );
  AND2X1_RVT U3163 ( .A1(n1910), .A2(N1129), .Y(\sub_381/carry[2] ) );
  XOR2X1_RVT U3164 ( .A1(N1188), .A2(N1129), .Y(N1595) );
  XNOR2X1_RVT U3165 ( .A1(n1926), .A2(\sub_312/carry[9] ), .Y(N1318) );
  OR2X1_RVT U3166 ( .A1(n1528), .A2(\sub_312/carry[8] ), .Y(\sub_312/carry[9] ) );
  XNOR2X1_RVT U3167 ( .A1(\sub_312/carry[8] ), .A2(n1923), .Y(N1317) );
  OR2X1_RVT U3168 ( .A1(n1922), .A2(\sub_312/carry[7] ), .Y(\sub_312/carry[8] ) );
  XNOR2X1_RVT U3169 ( .A1(\sub_312/carry[7] ), .A2(n1525), .Y(N1316) );
  OR2X1_RVT U3170 ( .A1(n1920), .A2(\sub_312/carry[6] ), .Y(\sub_312/carry[7] ) );
  XNOR2X1_RVT U3171 ( .A1(\sub_312/carry[6] ), .A2(n1527), .Y(N1315) );
  OR2X1_RVT U3172 ( .A1(n1918), .A2(n1914), .Y(\sub_312/carry[6] ) );
  XNOR2X1_RVT U3173 ( .A1(n1913), .A2(n1526), .Y(N1314) );
  XNOR2X1_RVT U3174 ( .A1(n1926), .A2(\sub_376/carry[9] ), .Y(N1593) );
  OR2X1_RVT U3175 ( .A1(n1528), .A2(\sub_376/carry[8] ), .Y(\sub_376/carry[9] ) );
  XNOR2X1_RVT U3176 ( .A1(\sub_376/carry[8] ), .A2(n1923), .Y(N1592) );
  OR2X1_RVT U3177 ( .A1(n1922), .A2(\sub_376/carry[7] ), .Y(\sub_376/carry[8] ) );
  XNOR2X1_RVT U3178 ( .A1(\sub_376/carry[7] ), .A2(n1525), .Y(N1591) );
  OR2X1_RVT U3179 ( .A1(n1920), .A2(\sub_376/carry[6] ), .Y(\sub_376/carry[7] ) );
  XNOR2X1_RVT U3180 ( .A1(\sub_376/carry[6] ), .A2(n1527), .Y(N1590) );
  OR2X1_RVT U3181 ( .A1(n1918), .A2(\sub_376/carry[5] ), .Y(\sub_376/carry[6] ) );
  XNOR2X1_RVT U3182 ( .A1(\sub_376/carry[5] ), .A2(n1526), .Y(N1589) );
  OR2X1_RVT U3183 ( .A1(n1915), .A2(n1903), .Y(\sub_376/carry[5] ) );
  XNOR2X1_RVT U3184 ( .A1(n1902), .A2(n1913), .Y(N1588) );
  XOR2X1_RVT U3185 ( .A1(n1528), .A2(\add_489/carry[8] ), .Y(N2053) );
  AND2X1_RVT U3186 ( .A1(n1922), .A2(\add_489/carry[7] ), .Y(
        \add_489/carry[8] ) );
  XOR2X1_RVT U3187 ( .A1(n1525), .A2(\add_489/carry[7] ), .Y(N2052) );
  OR2X1_RVT U3188 ( .A1(n1920), .A2(\add_489/carry[6] ), .Y(\add_489/carry[7] ) );
  XNOR2X1_RVT U3189 ( .A1(\add_489/carry[6] ), .A2(n1527), .Y(N2051) );
  OR2X1_RVT U3190 ( .A1(n1918), .A2(\add_489/carry[5] ), .Y(\add_489/carry[6] ) );
  XNOR2X1_RVT U3191 ( .A1(\add_489/carry[5] ), .A2(n1526), .Y(N2050) );
  OR2X1_RVT U3192 ( .A1(n1915), .A2(\add_489/carry[4] ), .Y(\add_489/carry[5] ) );
  XNOR2X1_RVT U3193 ( .A1(\add_489/carry[4] ), .A2(n1913), .Y(N2049) );
  OR2X1_RVT U3194 ( .A1(n1903), .A2(\add_489/carry[3] ), .Y(\add_489/carry[4] ) );
  XNOR2X1_RVT U3195 ( .A1(\add_489/carry[3] ), .A2(n1902), .Y(N2048) );
  OR2X1_RVT U3196 ( .A1(n1907), .A2(n1909), .Y(\add_489/carry[3] ) );
  XNOR2X1_RVT U3197 ( .A1(n1909), .A2(n1906), .Y(N2047) );
  XOR2X1_RVT U3198 ( .A1(n1927), .A2(\add_480/carry[9] ), .Y(N2044) );
  AND2X1_RVT U3199 ( .A1(n1924), .A2(\add_480/carry[8] ), .Y(
        \add_480/carry[9] ) );
  XOR2X1_RVT U3200 ( .A1(n1528), .A2(\add_480/carry[8] ), .Y(N2043) );
  AND2X1_RVT U3201 ( .A1(n1922), .A2(\add_480/carry[7] ), .Y(
        \add_480/carry[8] ) );
  XOR2X1_RVT U3202 ( .A1(n1525), .A2(\add_480/carry[7] ), .Y(N2042) );
  OR2X1_RVT U3203 ( .A1(n1920), .A2(\add_480/carry[6] ), .Y(\add_480/carry[7] ) );
  XNOR2X1_RVT U3204 ( .A1(\add_480/carry[6] ), .A2(n1527), .Y(N2041) );
  OR2X1_RVT U3205 ( .A1(n1918), .A2(\add_480/carry[5] ), .Y(\add_480/carry[6] ) );
  XNOR2X1_RVT U3206 ( .A1(\add_480/carry[5] ), .A2(n1526), .Y(N2040) );
  OR2X1_RVT U3207 ( .A1(n1915), .A2(\add_480/carry[4] ), .Y(\add_480/carry[5] ) );
  XNOR2X1_RVT U3208 ( .A1(\add_480/carry[4] ), .A2(n1913), .Y(N2039) );
  OR2X1_RVT U3209 ( .A1(n1903), .A2(\add_480/carry[3] ), .Y(\add_480/carry[4] ) );
  XNOR2X1_RVT U3210 ( .A1(\add_480/carry[3] ), .A2(n1902), .Y(N2038) );
  OR2X1_RVT U3211 ( .A1(n1907), .A2(\add_480/carry[2] ), .Y(\add_480/carry[3] ) );
  XNOR2X1_RVT U3212 ( .A1(\add_480/carry[2] ), .A2(n1906), .Y(N2037) );
  OR2X1_RVT U3213 ( .A1(n1909), .A2(N1129), .Y(\add_480/carry[2] ) );
  XNOR2X1_RVT U3214 ( .A1(N1129), .A2(n1909), .Y(N2036) );
  XNOR2X1_RVT U3215 ( .A1(n1926), .A2(\sub_458/carry[9] ), .Y(N1965) );
  OR2X1_RVT U3216 ( .A1(n1924), .A2(\sub_458/carry[8] ), .Y(\sub_458/carry[9] ) );
  XNOR2X1_RVT U3217 ( .A1(\sub_458/carry[8] ), .A2(n1923), .Y(N1964) );
  OR2X1_RVT U3218 ( .A1(n1922), .A2(\sub_458/carry[7] ), .Y(\sub_458/carry[8] ) );
  XNOR2X1_RVT U3219 ( .A1(\sub_458/carry[7] ), .A2(n1525), .Y(N1963) );
  AND2X1_RVT U3220 ( .A1(n1920), .A2(\sub_458/carry[6] ), .Y(
        \sub_458/carry[7] ) );
  XOR2X1_RVT U3221 ( .A1(n1527), .A2(\sub_458/carry[6] ), .Y(N1962) );
  AND2X1_RVT U3222 ( .A1(n1918), .A2(\sub_458/carry[5] ), .Y(
        \sub_458/carry[6] ) );
  XOR2X1_RVT U3223 ( .A1(n1526), .A2(\sub_458/carry[5] ), .Y(N1961) );
  AND2X1_RVT U3224 ( .A1(n1916), .A2(\sub_458/carry[4] ), .Y(
        \sub_458/carry[5] ) );
  XOR2X1_RVT U3225 ( .A1(n1914), .A2(\sub_458/carry[4] ), .Y(N1960) );
  AND2X1_RVT U3226 ( .A1(n1904), .A2(\sub_458/carry[3] ), .Y(
        \sub_458/carry[4] ) );
  XOR2X1_RVT U3227 ( .A1(n1903), .A2(\sub_458/carry[3] ), .Y(N1959) );
  AND2X1_RVT U3228 ( .A1(n1908), .A2(n1910), .Y(\sub_458/carry[3] ) );
  XOR2X1_RVT U3229 ( .A1(n1907), .A2(n1909), .Y(N1958) );
  OR2X1_RVT U3230 ( .A1(n1910), .A2(n1911), .Y(n2327) );
  AO21X1_RVT U3231 ( .A1(n1910), .A2(N1129), .A3(n2335), .Y(N1820) );
  OR2X1_RVT U3232 ( .A1(n2327), .A2(n1907), .Y(n2328) );
  AO21X1_RVT U3233 ( .A1(n1908), .A2(n2327), .A3(n2336), .Y(N1821) );
  OR2X1_RVT U3234 ( .A1(n2328), .A2(n1903), .Y(n2329) );
  AO21X1_RVT U3235 ( .A1(n1905), .A2(n2328), .A3(n2337), .Y(N1822) );
  OR2X1_RVT U3236 ( .A1(n2329), .A2(n1914), .Y(n2330) );
  AO21X1_RVT U3237 ( .A1(n1916), .A2(n2329), .A3(n2338), .Y(N1823) );
  OR2X1_RVT U3238 ( .A1(n2330), .A2(n1526), .Y(n2331) );
  AO21X1_RVT U3239 ( .A1(n1918), .A2(n2330), .A3(n2339), .Y(N1824) );
  OR2X1_RVT U3240 ( .A1(n2331), .A2(n1527), .Y(n2332) );
  AO21X1_RVT U3241 ( .A1(n1920), .A2(n2331), .A3(n2340), .Y(N1825) );
  NOR2X0_RVT U3242 ( .A1(n2332), .A2(n1525), .Y(n2333) );
  AO21X1_RVT U3243 ( .A1(n1922), .A2(n2332), .A3(n2333), .Y(N1826) );
  XNOR2X1_RVT U3244 ( .A1(n1594), .A2(n2333), .Y(N1827) );
  NAND2X0_RVT U3245 ( .A1(n2333), .A2(n1594), .Y(n2334) );
  XNOR2X1_RVT U3246 ( .A1(n2334), .A2(n1927), .Y(N1828) );
  NAND2X0_RVT U3247 ( .A1(a_e[5]), .A2(n1537), .Y(n2363) );
  OR2X1_RVT U3248 ( .A1(n1261), .A2(b_e[4]), .Y(n2347) );
  NAND2X0_RVT U3249 ( .A1(a_e[3]), .A2(n1536), .Y(n2358) );
  OR2X1_RVT U3250 ( .A1(n1257), .A2(b_e[2]), .Y(n2344) );
  NAND2X0_RVT U3251 ( .A1(a_e[0]), .A2(n1539), .Y(n2341) );
  OR2X1_RVT U3252 ( .A1(n2341), .A2(n1255), .Y(n2342) );
  NAND2X0_RVT U3253 ( .A1(b_e[2]), .A2(n1257), .Y(n2355) );
  NAND2X0_RVT U3254 ( .A1(n2344), .A2(n2355), .Y(n2351) );
  AO221X1_RVT U3255 ( .A1(b_e[1]), .A2(n2342), .A3(n2341), .A4(n1255), .A5(
        n2351), .Y(n2343) );
  NAND3X0_RVT U3256 ( .A1(n2358), .A2(n2344), .A3(n2343), .Y(n2345) );
  OR2X1_RVT U3257 ( .A1(n1536), .A2(a_e[3]), .Y(n2354) );
  NAND2X0_RVT U3258 ( .A1(b_e[4]), .A2(n1261), .Y(n2361) );
  AND2X1_RVT U3259 ( .A1(n2347), .A2(n2361), .Y(n2357) );
  NAND3X0_RVT U3260 ( .A1(n2345), .A2(n2354), .A3(n2357), .Y(n2346) );
  NAND3X0_RVT U3261 ( .A1(n2363), .A2(n2347), .A3(n2346), .Y(n2348) );
  OR2X1_RVT U3262 ( .A1(n1537), .A2(a_e[5]), .Y(n2360) );
  AND2X1_RVT U3263 ( .A1(n2348), .A2(n2360), .Y(n2349) );
  XNOR2X1_RVT U3264 ( .A1(a_e[6]), .A2(b_e[6]), .Y(n2365) );
  AO22X1_RVT U3265 ( .A1(n2349), .A2(n2365), .A3(a_e[6]), .A4(n1535), .Y(n2350) );
  NAND2X0_RVT U3266 ( .A1(b_e[7]), .A2(n1267), .Y(n2367) );
  OR2X1_RVT U3267 ( .A1(n1267), .A2(b_e[7]), .Y(n2368) );
  AO21X1_RVT U3268 ( .A1(n2350), .A2(n2367), .A3(n2370), .Y(N95) );
  OR2X1_RVT U3269 ( .A1(n1539), .A2(a_e[0]), .Y(n2352) );
  OR2X1_RVT U3270 ( .A1(n2352), .A2(a_e[1]), .Y(n2353) );
  AO221X1_RVT U3271 ( .A1(n2353), .A2(n1538), .A3(a_e[1]), .A4(n2352), .A5(
        n2351), .Y(n2356) );
  NAND3X0_RVT U3272 ( .A1(n2356), .A2(n2355), .A3(n2354), .Y(n2359) );
  NAND3X0_RVT U3273 ( .A1(n2359), .A2(n2358), .A3(n2357), .Y(n2362) );
  NAND3X0_RVT U3274 ( .A1(n2362), .A2(n2361), .A3(n2360), .Y(n2364) );
  AND2X1_RVT U3275 ( .A1(n2364), .A2(n2363), .Y(n2366) );
  AO22X1_RVT U3276 ( .A1(n2366), .A2(n2365), .A3(b_e[6]), .A4(n1265), .Y(n2369) );
  AO21X1_RVT U3277 ( .A1(n2369), .A2(n2368), .A3(n2371), .Y(N94) );
  XNOR2X1_RVT U3278 ( .A1(tmp_b_e1[6]), .A2(tmp_a_e1[6]), .Y(n2375) );
  XNOR2X1_RVT U3279 ( .A1(tmp_b_e1[5]), .A2(tmp_a_e1[5]), .Y(n2374) );
  XNOR2X1_RVT U3280 ( .A1(tmp_b_e1[4]), .A2(tmp_a_e1[4]), .Y(n2373) );
  XNOR2X1_RVT U3281 ( .A1(tmp_b_e1[3]), .A2(tmp_a_e1[3]), .Y(n2372) );
  NAND4X0_RVT U3282 ( .A1(n2375), .A2(n2374), .A3(n2373), .A4(n2372), .Y(n2383) );
  XNOR2X1_RVT U3283 ( .A1(tmp_b_e1[2]), .A2(tmp_a_e1[2]), .Y(n2377) );
  XNOR2X1_RVT U3284 ( .A1(tmp_b_e1[7]), .A2(tmp_a_e1[7]), .Y(n2376) );
  NAND2X0_RVT U3285 ( .A1(n2377), .A2(n2376), .Y(n2382) );
  NOR2X0_RVT U3286 ( .A1(n2384), .A2(tmp_a_e1[0]), .Y(n2378) );
  OA22X1_RVT U3287 ( .A1(tmp_b_e1[1]), .A2(n2378), .A3(n2378), .A4(n2456), .Y(
        n2381) );
  AND2X1_RVT U3288 ( .A1(tmp_a_e1[0]), .A2(n2384), .Y(n2379) );
  OA22X1_RVT U3289 ( .A1(n2379), .A2(n2385), .A3(tmp_a_e1[1]), .A4(n2379), .Y(
        n2380) );
  NOR4X0_RVT U3290 ( .A1(n2383), .A2(n2382), .A3(n2381), .A4(n2380), .Y(N2131)
         );
  XNOR2X1_RVT U3291 ( .A1(tmp_b_m1[4]), .A2(tmp_a_m1[4]), .Y(n2394) );
  XNOR2X1_RVT U3292 ( .A1(tmp_b_m1[3]), .A2(tmp_a_m1[3]), .Y(n2393) );
  XNOR2X1_RVT U3293 ( .A1(tmp_b_m1[5]), .A2(tmp_a_m1[5]), .Y(n2392) );
  XOR2X1_RVT U3294 ( .A1(tmp_b_m1[2]), .A2(tmp_a_m1[2]), .Y(n2390) );
  NOR2X0_RVT U3295 ( .A1(n2463), .A2(tmp_b_m1[0]), .Y(n2386) );
  OA22X1_RVT U3296 ( .A1(n2386), .A2(n2420), .A3(tmp_a_m1[1]), .A4(n2386), .Y(
        n2389) );
  AND2X1_RVT U3297 ( .A1(tmp_b_m1[0]), .A2(n2463), .Y(n2387) );
  OA22X1_RVT U3298 ( .A1(tmp_b_m1[1]), .A2(n2387), .A3(n2387), .A4(n2419), .Y(
        n2388) );
  NOR3X0_RVT U3299 ( .A1(n2390), .A2(n2389), .A3(n2388), .Y(n2391) );
  NAND4X0_RVT U3300 ( .A1(n2394), .A2(n2393), .A3(n2392), .A4(n2391), .Y(n2418) );
  XNOR2X1_RVT U3301 ( .A1(tmp_b_m1[10]), .A2(tmp_a_m1[10]), .Y(n2401) );
  XNOR2X1_RVT U3302 ( .A1(tmp_b_m1[9]), .A2(tmp_a_m1[9]), .Y(n2400) );
  XNOR2X1_RVT U3303 ( .A1(tmp_b_m1[11]), .A2(tmp_a_m1[11]), .Y(n2399) );
  XNOR2X1_RVT U3304 ( .A1(tmp_b_m1[7]), .A2(tmp_a_m1[7]), .Y(n2397) );
  XNOR2X1_RVT U3305 ( .A1(tmp_b_m1[6]), .A2(tmp_a_m1[6]), .Y(n2396) );
  XNOR2X1_RVT U3306 ( .A1(tmp_b_m1[8]), .A2(tmp_a_m1[8]), .Y(n2395) );
  AND3X1_RVT U3307 ( .A1(n2397), .A2(n2396), .A3(n2395), .Y(n2398) );
  NAND4X0_RVT U3308 ( .A1(n2401), .A2(n2400), .A3(n2399), .A4(n2398), .Y(n2417) );
  XNOR2X1_RVT U3309 ( .A1(tmp_b_m1[16]), .A2(tmp_a_m1[16]), .Y(n2408) );
  XNOR2X1_RVT U3310 ( .A1(tmp_b_m1[15]), .A2(tmp_a_m1[15]), .Y(n2407) );
  XNOR2X1_RVT U3311 ( .A1(tmp_b_m1[17]), .A2(tmp_a_m1[17]), .Y(n2406) );
  XNOR2X1_RVT U3312 ( .A1(tmp_b_m1[13]), .A2(tmp_a_m1[13]), .Y(n2404) );
  XNOR2X1_RVT U3313 ( .A1(tmp_b_m1[12]), .A2(tmp_a_m1[12]), .Y(n2403) );
  XNOR2X1_RVT U3314 ( .A1(tmp_b_m1[14]), .A2(tmp_a_m1[14]), .Y(n2402) );
  AND3X1_RVT U3315 ( .A1(n2404), .A2(n2403), .A3(n2402), .Y(n2405) );
  NAND4X0_RVT U3316 ( .A1(n2408), .A2(n2407), .A3(n2406), .A4(n2405), .Y(n2416) );
  XNOR2X1_RVT U3317 ( .A1(tmp_b_m1[19]), .A2(tmp_a_m1[19]), .Y(n2414) );
  XNOR2X1_RVT U3318 ( .A1(tmp_b_m1[18]), .A2(tmp_a_m1[18]), .Y(n2413) );
  XNOR2X1_RVT U3319 ( .A1(tmp_b_m1[20]), .A2(tmp_a_m1[20]), .Y(n2412) );
  XNOR2X1_RVT U3320 ( .A1(tmp_b_m1[22]), .A2(tmp_a_m1[22]), .Y(n2410) );
  XNOR2X1_RVT U3321 ( .A1(tmp_b_m1[21]), .A2(tmp_a_m1[21]), .Y(n2409) );
  AND2X1_RVT U3322 ( .A1(n2410), .A2(n2409), .Y(n2411) );
  NAND4X0_RVT U3323 ( .A1(n2414), .A2(n2413), .A3(n2412), .A4(n2411), .Y(n2415) );
  NOR4X0_RVT U3324 ( .A1(n2418), .A2(n2417), .A3(n2416), .A4(n2415), .Y(N2132)
         );
  AND4X1_RVT U3325 ( .A1(tmp_e1[4]), .A2(tmp_e1[3]), .A3(tmp_e1[7]), .A4(
        tmp_e1[6]), .Y(n2421) );
  OR3X1_RVT U3326 ( .A1(N2211), .A2(N2210), .A3(N2209), .Y(n2422) );
  NOR4X0_RVT U3327 ( .A1(n2422), .A2(N2206), .A3(N2208), .A4(N2207), .Y(n2429)
         );
  OR3X1_RVT U3328 ( .A1(N2217), .A2(N2216), .A3(N2215), .Y(n2423) );
  NOR4X0_RVT U3329 ( .A1(n2423), .A2(N2212), .A3(N2214), .A4(N2213), .Y(n2428)
         );
  OR3X1_RVT U3330 ( .A1(N2223), .A2(N2222), .A3(N2221), .Y(n2424) );
  NOR4X0_RVT U3331 ( .A1(n2424), .A2(N2218), .A3(N2220), .A4(N2219), .Y(n2427)
         );
  OR3X1_RVT U3332 ( .A1(N2450), .A2(N2228), .A3(N2227), .Y(n2425) );
  NOR4X0_RVT U3333 ( .A1(n2425), .A2(N2224), .A3(N2226), .A4(N2225), .Y(n2426)
         );
  NAND4X0_RVT U3334 ( .A1(n2429), .A2(n2428), .A3(n2427), .A4(n2426), .Y(N2230) );
  NOR4X0_RVT U3335 ( .A1(tmp_e1[3]), .A2(tmp_e1[2]), .A3(tmp_e1[1]), .A4(
        tmp_e1[0]), .Y(n2432) );
  OR2X1_RVT U3336 ( .A1(tmp_e1[8]), .A2(tmp_e1[7]), .Y(n2430) );
  NOR4X0_RVT U3337 ( .A1(tmp_e1[6]), .A2(n2430), .A3(tmp_e1[5]), .A4(tmp_e1[4]), .Y(n2431) );
  AO21X1_RVT U3338 ( .A1(n2432), .A2(n2431), .A3(tmp_e1[9]), .Y(N2119) );
  NAND4X0_RVT U3339 ( .A1(tmp_e1[1]), .A2(tmp_e1[0]), .A3(tmp_e1[5]), .A4(
        tmp_e1[2]), .Y(n2434) );
  NAND4X0_RVT U3340 ( .A1(tmp_e1[4]), .A2(tmp_e1[3]), .A3(tmp_e1[7]), .A4(
        tmp_e1[6]), .Y(n2433) );
  NOR2X0_RVT U3341 ( .A1(n2434), .A2(n2433), .Y(n2435) );
  OA21X1_RVT U3342 ( .A1(tmp_e1[8]), .A2(n2435), .A3(n1784), .Y(N2118) );
endmodule
