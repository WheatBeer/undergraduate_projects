`timescale 1ns/100ps

module test;
    reg clk;
    reg rst;
    reg [31:0] a;
    reg [31:0] b;
    reg [1:0] sel;
    wire err;
    wire overflow;
    wire [31:0] y;

    fpu fpu_test(clk, rst, a, b, sel, err, overflow, y);

    always // clock generation
    begin
        #5 clk = ~clk;
    end

    initial
    begin
        clk <= 1;
        rst <= 0;
        a <= 0;
        b <= 0;
        sel <= 0;

/*************** sel = 0: add ***************/
// all exception case

        #9
        // y =  nan
        a <= 32'b0_11111111_00000000000000000000000;  // a =  inf
        b <= 32'b0_11111111_00000000000000000000000;  // b =  inf

        #10
        // y =  -nan
        a <= 32'b1_11111111_00000000000000000000000;  // a =  -inf
        b <= 32'b0_11111111_00000000000000000000000;  // b =  inf

        #10
        // y =  nan
        a <= 32'b0_11111111_10000000000000000000000;  // a =  nan
        b <= 32'b0_01111111_00000000000000000000000;  // b =  1.0

        #10
        sel <= 2'b00;
        // y =  0.00
        a <= 32'b0_00000000_00000000000000000000000;  // a =  0.0
        b <= 32'b0_00000000_00000000000000000000000;  // b =  0.0

        #10
        // y =  overflow, +inf
        a <= 32'b0_11111110_10100100001001000000000;  // a =  2.7923134E38(very large number)
        b <= 32'b0_11111110_11110100001001000000000;  // b =  3.3240046E38(very large number)

        #10
        // y =  overflow, -inf
        a <= 32'b1_11111110_10100100001001000000000;  // a =  -2.7923134E38(very large number)
        b <= 32'b1_11111110_11110100001001000000000;  // b =  -3.3240046E38(very large number)

        #10
        // y =  underflow, -0
        a <= 32'b0_00000000_00000000000000000000010;  // a =  2.8E-45(very small number)
        b <= 32'b1_00000000_00000000000000000000011;  // b =  -4.2E-45(very small number)

// all general case

        #10
        // y =  4.50
        a <= 32'b0_10000000_10000000000000000000000;  // a =  3.0
        b <= 32'b0_01111111_10000000000000000000000;  // b =  1.5

        #10
        // y =  6.0
        a <= 32'b0_10000000_10000000000000000000000;  // a =  3.0
        b <= 32'b0_10000000_10000000000000000000000;  // a =  3.0

        #10
        // y =  -1.20
        a <= 32'b0_01111101_00110100001110010101100;  // a =  0.301
        b <= 32'b1_01111111_10000000000000000000000;  // b =  -1.5

        #10
        // y =  -1411.40
        a <= 32'b1_10001001_01100000100000000000000;  // a =  -1410.0
        b <= 32'b1_01111111_01100110011001100110011;  // b =  -1.4

        #10
        // y =  1760
        a <= 32'b0_10001000_11111000000000000000000;  // a =  1008
        b <= 32'b0_10001000_01111000000000000000000;  // b =  752

        #10
        // y =  1056
        a <= 32'b0_10001000_00010000000000000000000;  // a =  544
        b <= 32'b0_10001000_00000000000000000000000;  // b =  512 

        #10
        // y =  2560
        a <= 32'b0_10001001_00000000000000000000000;  // a =  1024
        b <= 32'b0_10001010_10000000000000000000000;  // b =  1536
        
        #10
        // y =  131072.25
        a <= 32'b0_10001111_00000000000000000010000;  // a =  65536.125
        b <= 32'b0_10001111_00000000000000000010000;  // b =  65536.125
        
        
/*************** sel = 1: sub ***************/

// all exception case
        #10
        sel <= 2'b01;
        // y =  0.00
        a <= 32'b0_00000000_00000000000000000000000;  // a =  0.0
        b <= 32'b0_00000000_00000000000000000000000;  // b =  0.0

        #10
        // y =  inf
        a <= 32'b0_11111111_00000000000000000000000;  // a =  inf
        b <= 32'b0_11111111_00000000000000000000000;  // b =  inf

        #10
        // y =  -inf
        a <= 32'b1_11111111_00000000000000000000000;  // a =  -inf
        b <= 32'b0_11111111_00000000000000000000000;  // b =  inf

        #10
        // y =  nan
        a <= 32'b0_11111111_10000000000000000000000;  // a =  nan
        b <= 32'b0_01111111_00000000000000000000000;  // b =  1.0


        #10
        // y =  overflow, +inf
        a <= 32'b0_11111110_10100100001001000000000;  // a =  2.7923134E38(very large number)
        b <= 32'b1_11111110_11110100001001000000000;  // b = -3.3240046E38(very large number)

        #10
        // y =  overflow, -inf
        a <= 32'b1_11111110_10100100001001000000000;  // a =  -2.7923134E38(very large number)
        b <= 32'b0_11111110_11110100001001000000000;  // b =  3.3240046E38(very large number)

        #10
        // y =  underflow, +0
        a <= 32'b1_00000000_00000000000000000000010;  // a =  -2.8E-45(very small number)
        b <= 32'b1_00000000_00000000000000000000011;  // b =  -4.2E-45(very small number)


// all general case

        #10
        // y =  -0.11
        a <= 32'b0_01111111_01010100011110101110001;  // a =  1.33
        b <= 32'b0_01111111_01110000101000111101100;  // b =  1.44
        
        #10
        // y =  -2.77
        a <= 32'b1_01111111_01010100011110101110001;  // a =  -1.33
        b <= 32'b0_01111111_01110000101000111101100;  // b =  1.44

        #10
        // y =  2.67
        a <= 32'b0_01111101_01010001111010111000011;  // a =  0.33
        b <= 32'b1_10000000_00101011100001010001111;  // b =  -2.34

        #10
        // y =  2.01
        a <= 32'b1_01111101_01010001111010111000011;  // a =  -0.33
        b <= 32'b1_10000000_00101011100001010001111;  // b =  -2.34

        #10
        // y =  0
        a <= 32'b0_10000000_10000000000000000000000;  // a =  3.0
        b <= 32'b0_10000000_10000000000000000000000;  // a =  3.0
        
        #10
        a <= 32'b1_10001000_11111000000000000000000;  // a =  -1008
        b <= 32'b1_10001000_01111000000000000000000;  // b =  -752

        #10
        a <= 32'b1_10001000_00010000000000000000000;  // a =  -544
        b <= 32'b1_10001000_00000000000000000000000;  // b =  -512

        #10
        // y =  1024.250
        a <= 32'b0_10001000_00000000000100000000000;  // a =  512.125
        b <= 32'b1_10001000_00000000000100000000000;  // b =  -512.125
        
/*************** sel = 2: mul ***************/

// all exception case
        #10
        sel <= 2'b10;
        // y = NaN
        a <= 32'b0_11111111_00000000000000000000001; // a = NaN
        b <= 32'b0_01111011_10011001100110011001101; // b = 0.1

        #10
        // y = -inf
        a <= 32'b0_11111111_00000000000000000000000; // a = +inf
        b <= 32'b1_01111011_10011001100110011001101; // b = -0.1
        
        #10
        // y = NaN
        a <= 32'b1_11111111_00000000000000000000000; // a = -inf
        b <= 32'b0_00000000_00000000000000000000000; // b = +0

        #10
        // y = overflow, -inf
        a <= 32'b1_11111000_10101000000000000000000; // a = -4.4030677E36
        b <= 32'b0_11110110_10000000000000000000000; // b = 9.96921E35

        #10
        // y = underflow, -0
        a <= 32'b0_00000110_10000000000000000000000; // a = 5.642373E-37
        b <= 32'b1_00000011_11000000000000000000000; // b = -8.2284605E-38


        #10
        // y = overflow, inf
        a <= 32'b0_11111110_01000000000000000000000; // a is almost inf
        b <= 32'b0_10000010_01100011001100110011010; // b = 11.11

        #10
        // y = underflow, +0
        a <= 32'b0_00000001_00000000000000000000010;  // a is almost zero
        b <= 32'b0_00000001_00000000000000000000010;  // b is almost zero

// all general case

        #10
        // y =  4.50
        a <= 32'b0_10000000_10000000000000000000000;  // a =  3.0
        b <= 32'b0_01111111_10000000000000000000000;  // b =  1.5


        #10
        // y = -0, normal number * zero
        a <= 32'b0_01111011_10011001100110011001101; // a = 0.1
        b <= 32'b1_00000000_00000000000000000000000; // b = -0

        #10
        // y = 11.0
        a <= 32'b0_10000000_00011001100110011001101; // a = 2.2
        b <= 32'b0_10000001_01000000000000000000000; // b = 5
        
        #10
        // y = 0.4
        a <= 32'b0_10000000_00000000000000000000000; // a = 2.0
        b <= 32'b0_01111100_10011001100110011001101; // b = 0.2


        
/*************** sel = 3: div ***************/
// all exception case
        #10
        sel <= 2'b11;
        // y =  nan
        a <= 32'b0_11111111_10000000000000000000000;  // a =  nan
        b <= 32'b0_11111111_10000000000000000000000;  // b =  nan

        #10
        // y =  inf
        a <= 32'b0_00000000_00000000000000000000000;  // a =  +0
        b <= 32'b0_00000000_00000000000000000000000;  // b =  +0

        #10
        // y =  divide by zero
        a <= 32'b0_01111011_10011001100110011001101;  // a =  0.1
        b <= 32'b0_00000000_00000000000000000000000;  // b =  +0


        #10
        // y =  nan
        a <= 32'b0_01111011_10011001100110011001101;  // a =  0.1
        b <= 32'b0_11111111_10000000000000000000000;  // b =  nan

        #10
        // y = +inf
        a <= 32'b0_11111110_01000000000000000000000;  // a is almost inf
        b <= 32'b0_00000000_00000000000000000000101;  // b is almost zero



        #10
        // y = +0
        a <= 32'b0_00000000_00000000000000000000010;  // a is almost zero
        b <= 32'b0_11111110_01000000000000000000000;  // b is almost inf


// all general case

        #10
        // y =  -3.00
        a <= 32'b1_01111101_00110011001100110011010;  // a =  -0.3
        b <= 32'b0_01111011_10011001100110011001101;  // b =  0.1

        #10
        // y = -1    a=b
        a <= 32'b0_10000010_00000000000000000000000; // a = 8
        b <= 32'b1_10000010_00000000000000000000000; // b = -8

        #10
        // y = 0.5  a_e<b_e, tmp's msb=1
        a <= 32'b1_10000001_00000000000000000000000; // a = -4
        b <= 32'b1_10000010_00000000000000000000000; // b = -8
        
        #10
        // y = 0.71x a_m<b_m, tmp's msb=0
        a <= 32'b0_10000001_01000000000000000000000; // a = 5
        b <= 32'b0_10000001_11000000000000000000000; // b = 7
        
        #10
        // y = 0.333  a<b, tmp's msb=0
        a <= 32'b0_10000000_00000000000000000000000; // a = 2
        b <= 32'b0_10000001_10000000000000000000000; // b = 6

        #10
        // y = 3  a>b, tmp's msb=1
        a <= 32'b0_10000000_10000000000000000000000; // a = 3
        b <= 32'b0_01111111_00000000000000000000000; // b = 1
    end
endmodule
